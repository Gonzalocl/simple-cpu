//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "ETC.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
supply0 w43;    //: /sn:0 {0}(-82,-21)(-103,-21){1}
//: {2}(-105,-23)(-105,-30){3}
//: {4}(-103,-32)(-93,-32)(-93,-31)(-82,-31){5}
//: {6}(-105,-34)(-105,-60){7}
//: {8}(-103,-62)(-93,-62)(-93,-61)(-82,-61){9}
//: {10}(-105,-64)(-105,-71)(-82,-71){11}
//: {12}(-107,-62)(-117,-62)(-117,-51)(-82,-51){13}
//: {14}(-107,-32)(-117,-32)(-117,-41)(-82,-41){15}
//: {16}(-105,-19)(-105,-12){17}
wire w6;    //: /sn:0 {0}(421,233)(421,218){1}
wire [31:0] w32;    //: /sn:0 {0}(#:-348,299)(-358,299)(-358,766)(667,766)(667,319){1}
//: {2}(669,317)(766,317)(766,340)(#:779,340){3}
//: {4}(665,317)(#:630,317){5}
wire [31:0] w7;    //: /sn:0 {0}(#:207,-31)(#:240,-31){1}
wire [31:0] w93;    //: /sn:0 {0}(#:779,498)(764,498){1}
wire [31:0] w73;    //: /sn:0 {0}(#:360,30)(250,30){1}
//: {2}(248,28)(248,6)(-567,6)(-567,75){3}
//: {4}(-565,77)(#:-421,77){5}
//: {6}(-567,79)(-567,184)(#:-659,184){7}
//: {8}(248,32)(248,71)(#:778,71){9}
wire [31:0] w96;    //: /sn:0 {0}(#:1370,4)(1254,4)(1254,297){1}
//: {2}(1252,299)(#:1221,299){3}
//: {4}(1254,301)(1254,741)(263,741){5}
//: {6}(261,739)(261,367)(#:291,367){7}
//: {8}(259,741)(-510,741)(-510,97)(#:-421,97){9}
wire [2:0] w112;    //: /sn:0 {0}(#:209,223)(209,208){1}
wire [31:0] w99;    //: /sn:0 {0}(#:-421,183)(-436,183){1}
wire [31:0] w122;    //: /sn:0 {0}(#:1370,170)(1355,170){1}
wire [31:0] w16;    //: /sn:0 {0}(#:389,-31)(#:330,-31){1}
wire w14;    //: /sn:0 {0}(533,276)(518,276){1}
wire w15;    //: /sn:0 {0}(533,266)(518,266){1}
wire [4:0] w89;    //: /sn:0 {0}(#:-81,222)(22,222)(22,192)(76,192){1}
//: {2}(80,192)(148,192){3}
//: {4}(152,192)(318,192)(318,272)(#:359,272){5}
//: {6}(150,194)(150,240)(#:188,240){7}
//: {8}(#:78,190)(78,-26)(201,-26){9}
wire w19;    //: /sn:0 {0}(531,318)(516,318){1}
wire w4;    //: /sn:0 {0}(986,311)(1001,311){1}
wire [31:0] w81;    //: /sn:0 {0}(#:778,202)(763,202){1}
wire [3:0] w38;    //: /sn:0 {0}(616,-26)(528,-26)(#:528,35)(366,35){1}
wire [31:0] w106;    //: /sn:0 {0}(#:291,409)(276,409){1}
wire [31:0] w109;    //: /sn:0 {0}(#:291,498)(276,498){1}
wire [31:0] w129;    //: /sn:0 {0}(#:1370,-16)(1180,-16)(1180,111)(1048,111)(1048,273){1}
//: {2}(1050,275)(1109,275)(1109,290)(#:1122,290){3}
//: {4}(1046,275)(#:986,275){5}
wire [4:0] w114;    //: /sn:0 {0}(#:87,256)(#:188,256){1}
wire [31:0] w97;    //: /sn:0 {0}(#:-421,119)(-436,119){1}
wire w3;    //: /sn:0 {0}(986,293)(1077,293)(1077,92)(1136,92)(1136,-335)(-603,-335){1}
wire [2:0] w0;    //: /sn:0 {0}(#:917,261)(917,246){1}
wire [31:0] w37;    //: /sn:0 {0}(#:1412,54)(1683,54)(1683,-345)(-773,-345)(-773,175)(#:-758,175){1}
wire [31:0] w127;    //: /sn:0 {0}(#:622,-31)(1295,-31)(1295,26)(#:1370,26){1}
wire [4:0] w120;    //: /sn:0 {0}(#:188,367)(173,367){1}
wire [31:0] w34;    //: /sn:0 {0}(#:-265,286)(-242,286){1}
//: {2}(-240,284)(-240,208)(#:-213,208){3}
//: {4}(-240,288)(-240,369)(#:-205,369){5}
wire [31:0] w111;    //: /sn:0 {0}(#:291,553)(276,553){1}
wire [31:0] w76;    //: /sn:0 {0}(#:778,113)(763,113){1}
wire [31:0] w87;    //: /sn:0 {0}(750,360)(#:779,360){1}
wire [31:0] w102;    //: /sn:0 {0}(#:-421,263)(-436,263){1}
wire [31:0] w75;    //: /sn:0 {0}(#:632,265)(666,265)(666,91)(#:778,91){1}
wire w21;    //: /sn:0 {0}(-680,-316)(-695,-316){1}
wire [4:0] w119;    //: /sn:0 {0}(#:188,346)(173,346){1}
wire [31:0] w31;    //: /sn:0 {0}(#:-379,147)(-357,147)(-357,268)(#:-348,268){1}
wire [31:0] w100;    //: /sn:0 {0}(#:-421,208)(-436,208){1}
wire [31:0] w90;    //: /sn:0 {0}(595,683)(629,683)(#:629,408)(#:779,408){1}
wire [27:0] w28;    //: /sn:0 {0}(#:410,25)(366,25){1}
wire [3:0] w24;    //: /sn:0 {0}(#:497,-26)(395,-26){1}
wire [27:0] w20;    //: /sn:0 {0}(#:616,-36)(395,-36){1}
wire [31:0] w124;    //: /sn:0 {0}(#:1370,115)(1355,115){1}
wire w36;    //: /sn:0 {0}(-758,185)(-773,185){1}
wire w23;    //: /sn:0 {0}(-213,218)(-228,218){1}
wire [2:0] w41;    //: /sn:0 {0}(#:788,47)(788,32){1}
wire [31:0] w1;    //: /sn:0 {0}(#:820,141)(840,141)(840,281)(#:855,281){1}
wire [31:0] w108;    //: /sn:0 {0}(#:291,473)(276,473){1}
wire [31:0] w25;    //: /sn:0 {0}(#:-114,217)(#:-87,217){1}
wire [31:0] w126;    //: /sn:0 {0}(#:1370,52)(1355,52){1}
wire [31:0] w82;    //: /sn:0 {0}(#:778,229)(763,229){1}
wire [4:0] w116;    //: /sn:0 {0}(#:188,288)(173,288){1}
wire [31:0] w98;    //: /sn:0 {0}(#:-421,145)(-436,145){1}
wire [31:0] w125;    //: /sn:0 {0}(#:1370,90)(1355,90){1}
wire [2:0] w121;    //: /sn:0 {0}(#:1380,-40)(1380,-55){1}
wire [4:0] w118;    //: /sn:0 {0}(#:188,328)(173,328){1}
wire w40;    //: /sn:0 {0}(1122,300)(1107,300){1}
wire w18;    //: /sn:0 {0}(531,328)(516,328){1}
wire [31:0] w92;    //: /sn:0 {0}(#:779,471)(764,471){1}
wire w35;    //: /sn:0 {0}(-758,195)(-866,195)(-866,-319)(-716,-319){1}
wire [4:0] w8;    //: /sn:0 {0}(#:201,-36)(91,-36)(91,140){1}
//: {2}(93,142)(346,142)(346,251)(#:359,251){3}
//: {4}(89,142)(3,142)(3,212)(#:-81,212){5}
wire [31:0] w91;    //: /sn:0 {0}(#:779,446)(764,446){1}
wire [2:0] w103;    //: /sn:0 {0}(#:301,343)(301,328){1}
wire w30;    //: /sn:0 {0}(-309,248)(-309,233){1}
wire [31:0] w101;    //: /sn:0 {0}(#:-421,235)(-436,235){1}
wire w22;    //: /sn:0 {0}(-213,228)(-228,228){1}
wire w17;    //: /sn:0 {0}(-695,-321)(-653,-321)(-653,-333)(-624,-333){1}
wire [31:0] w123;    //: /sn:0 {0}(#:1370,142)(1355,142){1}
wire [4:0] w117;    //: /sn:0 {0}(#:188,311)(173,311){1}
wire [2:0] w84;    //: /sn:0 {0}(#:-411,53)(-411,38){1}
wire [2:0] w85;    //: /sn:0 {0}(#:789,316)(789,301){1}
wire w11;    //: /sn:0 {0}(424,347)(424,362){1}
wire [31:0] w12;    //: /sn:0 {0}(#:489,306)(512,306)(512,308)(#:531,308){1}
wire [31:0] w2;    //: /sn:0 {0}(#:821,410)(840,410)(840,305)(#:855,305){1}
wire [4:0] w77;    //: /sn:0 {0}(#:111,266)(87,266){1}
wire [31:0] w105;    //: /sn:0 {0}(#:-106,378)(-82,378)(-82,448)(255,448)(255,387)(#:291,387){1}
wire [31:0] w110;    //: /sn:0 {0}(#:291,525)(276,525){1}
wire [4:0] w115;    //: /sn:0 {0}(#:188,272)(173,272){1}
wire [31:0] w83;    //: /sn:0 {0}(#:778,257)(763,257){1}
wire [31:0] w10;    //: /sn:0 {0}(#:333,437)(344,437)(344,319)(#:359,319){1}
wire [31:0] w78;    //: /sn:0 {0}(#:778,139)(763,139){1}
wire [31:0] w13;    //: /sn:0 {0}(#:489,271)(509,271)(509,256)(#:533,256){1}
wire [31:0] w88;    //: /sn:0 {0}(#:779,382)(759,382)(759,391)(471,391)(471,681){1}
//: {2}(473,683)(505,683){3}
//: {4}(469,683)(436,683){5}
wire [31:0] w94;    //: /sn:0 {0}(#:779,526)(764,526){1}
wire w27;    //: /sn:0 {0}(-205,379)(-220,379){1}
wire w33;    //: /sn:0 {0}(-308,330)(-308,345){1}
wire w5;    //: /sn:0 {0}(-588,-330)(-603,-330){1}
wire [5:0] w29;    //: /sn:0 {0}(#:-76,-46)(#:201,-46){1}
wire [31:0] w107;    //: /sn:0 {0}(#:291,435)(276,435){1}
wire [15:0] w80;    //: /sn:0 {0}(#:81,266)(60,266){1}
//: {2}(#:58,264)(58,-16)(201,-16){3}
//: {4}(58,268)(58,314)(-52,314){5}
//: {6}(-54,312)(-54,232)(-81,232){7}
//: {8}(#:-54,316)(-54,683)(337,683){9}
wire [5:0] w42;    //: /sn:0 {0}(#:-81,202)(-2,202)(-2,60){1}
wire [4:0] w9;    //: /sn:0 {0}(#:230,323)(247,323)(247,297)(#:359,297){1}
wire [31:0] w79;    //: /sn:0 {0}(#:778,177)(763,177){1}
wire [5:0] w55;    //: /sn:0 {0}(#:109,276)(87,276){1}
wire w39;    //: /sn:0 {0}(1122,310)(1107,310){1}
wire w26;    //: /sn:0 {0}(-205,389)(-220,389){1}
//: enddecls

  //: comment g8 @(-704,167) /sn:0
  //: /line:"PC"
  //: /end
  Reg32bits g4 (.Din(w34), .Reloj(w23), .W(w22), .Dout(w25));   //: @(-212, 198) /sz:(97, 40) /sn:0 /p:[ Li0>3 Li1>0 Li2>0 Ro0<0 ]
  assign {w38, w28} = w73; //: CONCAT g55  @(361,30) /sn:0 /R:2 /w:[ 1 1 0 ] /dr:0 /tp:0 /drp:0
  //: joint g37 (w8) @(91, 142) /w:[ 2 1 4 -1 ]
  assign {w114, w77, w55} = w80; //: CONCAT g51  @(82,266) /sn:0 /R:2 /w:[ 0 1 1 0 ] /dr:1 /tp:0 /drp:0
  Reg32bits g13 (.Din(w129), .Reloj(w40), .W(w39), .Dout(w96));   //: @(1123, 280) /sz:(97, 40) /sn:0 /p:[ Li0>3 Li1>0 Li2>0 Ro0<3 ]
  Reg32bits g3 (.Din(w12), .Reloj(w19), .W(w18), .Dout(w32));   //: @(532, 298) /sz:(97, 40) /sn:0 /p:[ Li0>1 Li1>0 Li2>0 Ro0<5 ]
  //: comment g34 @(334,452) /sn:0
  //: /line:"0. Suma... (4a)"
  //: /line:"1. lw (5)"
  //: /end
  Reg32bits g2 (.Din(w13), .Reloj(w15), .W(w14), .Dout(w75));   //: @(534, 246) /sz:(97, 40) /sn:0 /p:[ Li0>1 Li1>0 Li2>0 Ro0<0 ]
  Banco32Reg g1 (.W(w6), .Esc(w10), .RegEsc(w9), .RegLeer1(w8), .RegLeer2(w89), .Reloj(w11), .Leer1(w13), .Leer2(w12));   //: @(360, 234) /sz:(128, 112) /sn:0 /p:[ Ti0>0 Li0>1 Li1>1 Li2>3 Li3>5 Bi0>0 Ro0<0 Ro1<0 ]
  //: joint g16 (w80) @(-54, 314) /w:[ 5 6 -1 8 ]
  //: comment g11 @(588,248) /sn:0
  //: /line:"A"
  //: /end
  assign {w42, w8, w89, w80} = w25; //: CONCAT g50  @(-86,217) /sn:0 /R:2 /w:[ 0 5 0 7 1 ] /dr:1 /tp:0 /drp:0
  //: comment g10 @(-189,361) /sn:0
  //: /line:"Dato memoria"
  //: /end
  //: comment g28 @(825,415) /sn:0
  //: /line:"0. Suma... (3a), beq (3c)"
  //: /line:"1. Incrementa el PC en 4 (1)"
  //: /line:"2. lw y sw (3b)"
  //: /line:"3. Decodificacion (2)"
  //: /end
  //: joint g19 (w80) @(58, 266) /w:[ 1 2 -1 4 ]
  n4 g27 (.Sa(w87));   //: @(709, 340) /sz:(40, 40) /sn:0 /p:[ Ro0<0 ]
  Extensor16a32 g32 (.E(w80), .Sa(w88));   //: @(338, 667) /sz:(97, 40) /sn:0 /p:[ Li0>9 Ro0<5 ]
  assign {w24, w20} = w16; //: CONCAT g38  @(390,-31) /sn:0 /R:2 /w:[ 1 1 0 ] /dr:0 /tp:0 /drp:0
  Memoria g6 (.W(w30), .Esc(w32), .Direc(w31), .Reloj(w33), .Leer(w34));   //: @(-347, 249) /sz:(81, 80) /sn:0 /p:[ Ti0>0 Li0>0 Li1>1 Bi0>0 Ro0<0 ]
  //: comment g57 @(5,501) /sn:0
  //: /line:"Gonzalo Caparr�s L�iz"
  //: /end
  assign w127 = {w38, w20}; //: CONCAT g53  @(621,-31) /sn:0 /w:[ 0 0 0 ] /dr:1 /tp:0 /drp:1
  //: comment g9 @(-192,197) /sn:0
  //: /line:"Instruccion"
  //: /end
  Reg32bits g7 (.Din(w37), .Reloj(w36), .W(w35), .Dout(w73));   //: @(-757, 165) /sz:(97, 40) /sn:0 /p:[ Li0>1 Li1>0 Li2>0 Ro0<7 ]
  //: joint g15 (w89) @(150, 192) /w:[ 4 -1 3 6 ]
  Mux3x32 g20 (.C(w41), .E7(w83), .E6(w82), .E5(w81), .E4(w79), .E3(w78), .E2(w76), .E1(w75), .E0(w73), .Sa(w1));   //: @(779, 48) /sz:(40, 234) /sn:0 /p:[ Ti0>0 Li0>0 Li1>0 Li2>0 Li3>0 Li4>0 Li5>0 Li6>1 Li7>9 Ro0<0 ]
  //: joint g31 (w129) @(1048, 275) /w:[ 2 1 4 -1 ]
  assign w29 = {w43, w43, w43, w43, w43, w43}; //: CONCAT g39  @(-77,-46) /sn:0 /w:[ 0 11 9 13 15 5 0 ] /dr:0 /tp:0 /drp:1
  //: comment g43 @(-375,53) /sn:0
  //: /line:"0. Direccion del PC (1)"
  //: /line:"1. lw (4b), sw (4c)"
  //: /end
  _GGAND2 #(6) g48 (.I0(w5), .I1(w3), .Z(w17));   //: @(-614,-333) /sn:0 /R:2 /w:[ 1 1 1 ]
  Desplazador2 g17 (.E(w7), .Sa(w16));   //: @(241, -47) /sz:(88, 40) /sn:0 /p:[ Li0>1 Ro0<1 ]
  Mux3x32 g25 (.C(w121), .E0(w129), .E1(w96), .E2(w127), .E3(w126), .E4(w125), .E5(w124), .E6(w123), .E7(w122), .Sa(w37));   //: @(1371, -39) /sz:(40, 234) /sn:0 /p:[ Ti0>0 Li0>0 Li1>0 Li2>1 Li3>0 Li4>0 Li5>0 Li6>0 Li7>0 Ro0<0 ]
  //: comment g29 @(824,50) /sn:0
  //: /line:"0. Incrementa el PC en 4 (1), Decodificacion (2)"
  //: /line:"1. Suma... (3a), lw y sw (3b), beq (3c)"
  //: /end
  //: joint g52 (w43) @(-105, -21) /w:[ 1 2 -1 16 ]
  //: joint g42 (w88) @(471, 683) /w:[ 2 1 4 -1 ]
  //: joint g56 (w73) @(248, 30) /w:[ 1 2 -1 8 ]
  //: comment g14 @(1153,279) /sn:0
  //: /line:"ALUout"
  //: /end
  Reg32bits g5 (.Din(w34), .Reloj(w27), .W(w26), .Dout(w105));   //: @(-204, 359) /sz:(97, 40) /sn:0 /p:[ Li0>5 Li1>0 Li2>0 Ro0<0 ]
  //: joint g44 (w96) @(261, 741) /w:[ 5 6 8 -1 ]
  //: joint g47 (w96) @(1254, 299) /w:[ -1 1 2 4 ]
  //: joint g36 (w89) @(78, 192) /w:[ 2 8 1 -1 ]
  Mux3x5 g24 (.C(w112), .E7(w120), .E6(w119), .E5(w118), .E4(w117), .E3(w116), .E2(w115), .E1(w114), .E0(w89), .Sa(w9));   //: @(189, 224) /sz:(40, 160) /sn:0 /p:[ Ti0>0 Li0>0 Li1>0 Li2>0 Li3>0 Li4>0 Li5>0 Li6>1 Li7>7 Ro0<0 ]
  Mux3x32 g21 (.C(w85), .E7(w94), .E6(w93), .E5(w92), .E4(w91), .E3(w90), .E2(w88), .E1(w87), .E0(w32), .Sa(w2));   //: @(780, 317) /sz:(40, 234) /sn:0 /p:[ Ti0>0 Li0>0 Li1>0 Li2>0 Li3>0 Li4>1 Li5>0 Li6>1 Li7>3 Ro0<0 ]
  //: joint g41 (w43) @(-105, -62) /w:[ 8 10 12 7 ]
  Mux3x32 g23 (.C(w103), .E7(w111), .E6(w110), .E5(w109), .E4(w108), .E3(w107), .E2(w106), .E1(w105), .E0(w96), .Sa(w10));   //: @(292, 344) /sz:(40, 234) /sn:0 /p:[ Ti0>0 Li0>0 Li1>0 Li2>0 Li3>0 Li4>0 Li5>0 Li6>1 Li7>7 Ro0<0 ]
  //: joint g54 (w73) @(-567, 77) /w:[ 4 3 -1 6 ]
  //: GROUND g40 (w43) @(-105,-6) /sn:0 /w:[ 17 ]
  //: joint g45 (w43) @(-105, -32) /w:[ 4 6 14 3 ]
  //: joint g26 (w34) @(-240, 286) /w:[ -1 2 1 4 ]
  ALU g0 (.C(w0), .B(w2), .A(w1), .Sa(w129), .Overflow(w4), .Cero(w3));   //: @(856, 262) /sz:(129, 64) /sn:0 /p:[ Ti0>0 Li0>1 Li1>1 Ro0<5 Ro1<0 Ro2<0 ]
  Mux3x32 g22 (.C(w84), .E7(w102), .E6(w101), .E5(w100), .E4(w99), .E3(w98), .E2(w97), .E1(w96), .E0(w73), .Sa(w31));   //: @(-420, 54) /sz:(40, 234) /sn:0 /p:[ Ti0>0 Li0>0 Li1>0 Li2>0 Li3>0 Li4>0 Li5>0 Li6>9 Li7>5 Ro0<0 ]
  //: comment g35 @(165,385) /sn:0
  //: /line:"0. lw (5)"
  //: /line:"1. Suma... (4a)"
  //: /end
  //: joint g46 (w32) @(667, 317) /w:[ 2 -1 4 1 ]
  assign w7 = {w29, w8, w89, w80}; //: CONCAT g18  @(206,-31) /sn:0 /w:[ 0 1 0 9 3 ] /dr:0 /tp:0 /drp:1
  //: comment g12 @(583,300) /sn:0
  //: /line:"B"
  //: /end
  //: comment g30 @(1415,-38) /sn:0
  //: /line:"0. Incrementa el PC en 4 (1)"
  //: /line:"1. beq (3c)"
  //: /line:"2. Salto (3d)"
  //: /end
  Desplazador2 g33 (.E(w88), .Sa(w90));   //: @(506, 667) /sz:(88, 40) /sn:0 /p:[ Li0>3 Ro0<0 ]
  _GGOR2 #(6) g49 (.I0(w21), .I1(w17), .Z(w35));   //: @(-706,-319) /sn:0 /R:2 /w:[ 1 0 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin Mux5cableado
module Mux5cableado(E4, E8, E13, S5, S23, S26, E1, E11, E28, S18, E19, E6, S6, E7, S21, E20, E31, S7, S16, E17, E25, E29, S20, E14, S12, S15, E21, E23, S9, S8, S22, E0, E26, S14, S1, S17, S29, E3, S2, S19, E2, S27, E16, E10, E27, S0, E9, S25, E15, S11, S30, S10, S31, E5, S24, E24, S4, S28, E22, S3, S13, E12, E18, E30);
//: interface  /sz:(46, 1099) /bd:[ Li0>E31[31:0](1065/1099) Li1>E30[31:0](1032/1099) Li2>E29[31:0](999/1099) Li3>E28[31:0](965/1099) Li4>E27[31:0](932/1099) Li5>E26[31:0](899/1099) Li6>E25[31:0](865/1099) Li7>E24[31:0](832/1099) Li8>E23[31:0](799/1099) Li9>E22[31:0](765/1099) Li10>E21[31:0](732/1099) Li11>E20[31:0](699/1099) Li12>E19[31:0](666/1099) Li13>E18[31:0](632/1099) Li14>E17[31:0](599/1099) Li15>E16[31:0](566/1099) Li16>E15[31:0](532/1099) Li17>E14[31:0](499/1099) Li18>E13[31:0](466/1099) Li19>E12[31:0](432/1099) Li20>E11[31:0](399/1099) Li21>E10[31:0](366/1099) Li22>E9[31:0](333/1099) Li23>E8[31:0](299/1099) Li24>E7[31:0](266/1099) Li25>E6[31:0](233/1099) Li26>E5[31:0](199/1099) Li27>E4[31:0](166/1099) Li28>E3[31:0](133/1099) Li29>E2[31:0](99/1099) Li30>E1[31:0](66/1099) Li31>E0[31:0](33/1099) Ro0<S31[31:0](1065/1099) Ro1<S30[31:0](1032/1099) Ro2<S29[31:0](999/1099) Ro3<S28[31:0](965/1099) Ro4<S27[31:0](932/1099) Ro5<S26[31:0](899/1099) Ro6<S25[31:0](865/1099) Ro7<S24[31:0](832/1099) Ro8<S23[31:0](799/1099) Ro9<S22[31:0](765/1099) Ro10<S21[31:0](732/1099) Ro11<S20[31:0](699/1099) Ro12<S19[31:0](666/1099) Ro13<S18[31:0](632/1099) Ro14<S17[31:0](599/1099) Ro15<S16[31:0](566/1099) Ro16<S15[31:0](532/1099) Ro17<S14[31:0](499/1099) Ro18<S13[31:0](466/1099) Ro19<S12[31:0](432/1099) Ro20<S11[31:0](399/1099) Ro21<S10[31:0](366/1099) Ro22<S9[31:0](333/1099) Ro23<S8[31:0](299/1099) Ro24<S7[31:0](266/1099) Ro25<S6[31:0](233/1099) Ro26<S5[31:0](200/1099) Ro27<S4[31:0](166/1099) Ro28<S3[31:0](133/1099) Ro29<S2[31:0](99/1099) Ro30<S1[31:0](66/1099) Ro31<S0[31:0](33/1099) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output [31:0] S7;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E19;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S28;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [31:0] S13;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [31:0] S23;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [31:0] S1;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [31:0] S25;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E10;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S17;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E8;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S20;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E5;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
input [31:0] E26;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
input [31:0] E3;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
input [31:0] E15;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S29;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [31:0] S2;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E31;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
input [31:0] E14;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S0;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E27;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S10;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [31:0] S11;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [31:0] S8;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E20;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
input [31:0] E24;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
input [31:0] E21;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S16;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E28;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S5;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E13;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S30;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E7;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
input [31:0] E1;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
input [31:0] E30;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S12;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E2;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S26;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E4;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S31;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E25;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S19;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E29;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
input [31:0] E0;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S15;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E16;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S14;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [31:0] S3;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E17;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S24;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [31:0] S18;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [31:0] S27;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E22;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
input [31:0] E6;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
input [31:0] E12;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S4;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [31:0] S21;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E9;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
input [31:0] E18;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S6;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E23;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [31:0] S9;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [31:0] S22;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E11;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
wire w32;    //: /sn:0 {0}(1,1)(1,1){1}
wire w45;    //: /sn:0 {0}(1,1)(1,1){1}
wire w832;    //: /sn:0 {0}(1,1)(1,1){1}
wire w699;    //: /sn:0 {0}(1,1)(1,1){1}
wire w760;    //: /sn:0 {0}(1,1)(1,1){1}
wire w769;    //: /sn:0 {0}(1,1)(1,1){1}
wire w810;    //: /sn:0 {0}(1,1)(1,1){1}
wire w266;    //: /sn:0 {0}(1,1)(1,1){1}
wire w19;    //: /sn:0 {0}(1,1)(1,1){1}
wire w4;    //: /sn:0 {0}(1,1)(1,1){1}
wire w852;    //: /sn:0 {0}(1,1)(1,1){1}
wire w916;    //: /sn:0 {0}(1,1)(1,1){1}
wire w864;    //: /sn:0 {0}(1,1)(1,1){1}
wire w965;    //: /sn:0 {0}(1,1)(1,1){1}
wire w719;    //: /sn:0 {0}(1,1)(1,1){1}
wire w994;    //: /sn:0 {0}(1,1)(1,1){1}
wire w513;    //: /sn:0 {0}(1,1)(1,1){1}
wire w431;    //: /sn:0 {0}(1,1)(1,1){1}
wire w344;    //: /sn:0 {0}(1,1)(1,1){1}
wire w119;    //: /sn:0 {0}(1,1)(1,1){1}
wire w498;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1014;    //: /sn:0 {0}(1,1)(1,1){1}
wire w294;    //: /sn:0 {0}(1,1)(1,1){1}
wire w90;    //: /sn:0 {0}(1,1)(1,1){1}
wire w614;    //: /sn:0 {0}(1,1)(1,1){1}
wire w167;    //: /sn:0 {0}(1,1)(1,1){1}
wire w587;    //: /sn:0 {0}(1,1)(1,1){1}
wire w552;    //: /sn:0 {0}(1,1)(1,1){1}
wire w842;    //: /sn:0 {0}(1,1)(1,1){1}
wire w964;    //: /sn:0 {0}(1,1)(1,1){1}
wire w272;    //: /sn:0 {0}(1,1)(1,1){1}
wire w508;    //: /sn:0 {0}(1,1)(1,1){1}
wire w300;    //: /sn:0 {0}(1,1)(1,1){1}
wire w126;    //: /sn:0 {0}(1,1)(1,1){1}
wire w788;    //: /sn:0 {0}(1,1)(1,1){1}
wire w872;    //: /sn:0 {0}(1,1)(1,1){1}
wire w103;    //: /sn:0 {0}(1,1)(1,1){1}
wire w481;    //: /sn:0 {0}(1,1)(1,1){1}
wire w883;    //: /sn:0 {0}(1,1)(1,1){1}
wire w915;    //: /sn:0 {0}(1,1)(1,1){1}
wire w314;    //: /sn:0 {0}(1,1)(1,1){1}
wire w238;    //: /sn:0 {0}(1,1)(1,1){1}
wire w520;    //: /sn:0 {0}(1,1)(1,1){1}
wire w574;    //: /sn:0 {0}(1,1)(1,1){1}
wire w297;    //: /sn:0 {0}(1,1)(1,1){1}
wire w487;    //: /sn:0 {0}(1,1)(1,1){1}
wire w779;    //: /sn:0 {0}(1,1)(1,1){1}
wire w911;    //: /sn:0 {0}(1,1)(1,1){1}
wire w211;    //: /sn:0 {0}(1,1)(1,1){1}
wire w738;    //: /sn:0 {0}(1,1)(1,1){1}
wire w44;    //: /sn:0 {0}(1,1)(1,1){1}
wire w818;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1016;    //: /sn:0 {0}(1,1)(1,1){1}
wire w433;    //: /sn:0 {0}(1,1)(1,1){1}
wire w367;    //: /sn:0 {0}(1,1)(1,1){1}
wire w316;    //: /sn:0 {0}(1,1)(1,1){1}
wire w83;    //: /sn:0 {0}(1,1)(1,1){1}
wire w115;    //: /sn:0 {0}(1,1)(1,1){1}
wire w10;    //: /sn:0 {0}(1,1)(1,1){1}
wire w647;    //: /sn:0 {0}(1,1)(1,1){1}
wire w275;    //: /sn:0 {0}(1,1)(1,1){1}
wire w469;    //: /sn:0 {0}(1,1)(1,1){1}
wire w95;    //: /sn:0 {0}(1,1)(1,1){1}
wire w462;    //: /sn:0 {0}(1,1)(1,1){1}
wire w473;    //: /sn:0 {0}(1,1)(1,1){1}
wire w478;    //: /sn:0 {0}(1,1)(1,1){1}
wire w902;    //: /sn:0 {0}(1,1)(1,1){1}
wire w178;    //: /sn:0 {0}(1,1)(1,1){1}
wire w330;    //: /sn:0 {0}(1,1)(1,1){1}
wire w413;    //: /sn:0 {0}(1,1)(1,1){1}
wire w881;    //: /sn:0 {0}(1,1)(1,1){1}
wire w947;    //: /sn:0 {0}(1,1)(1,1){1}
wire w744;    //: /sn:0 {0}(1,1)(1,1){1}
wire w540;    //: /sn:0 {0}(1,1)(1,1){1}
wire w441;    //: /sn:0 {0}(1,1)(1,1){1}
wire w153;    //: /sn:0 {0}(1,1)(1,1){1}
wire w961;    //: /sn:0 {0}(1,1)(1,1){1}
wire w523;    //: /sn:0 {0}(1,1)(1,1){1}
wire w640;    //: /sn:0 {0}(1,1)(1,1){1}
wire w428;    //: /sn:0 {0}(1,1)(1,1){1}
wire w304;    //: /sn:0 {0}(1,1)(1,1){1}
wire w239;    //: /sn:0 {0}(1,1)(1,1){1}
wire w213;    //: /sn:0 {0}(1,1)(1,1){1}
wire w207;    //: /sn:0 {0}(1,1)(1,1){1}
wire w51;    //: /sn:0 {0}(1,1)(1,1){1}
wire w499;    //: /sn:0 {0}(1,1)(1,1){1}
wire w709;    //: /sn:0 {0}(1,1)(1,1){1}
wire w997;    //: /sn:0 {0}(1,1)(1,1){1}
wire w299;    //: /sn:0 {0}(1,1)(1,1){1}
wire w474;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1021;    //: /sn:0 {0}(1,1)(1,1){1}
wire w980;    //: /sn:0 {0}(1,1)(1,1){1}
wire w463;    //: /sn:0 {0}(1,1)(1,1){1}
wire w856;    //: /sn:0 {0}(1,1)(1,1){1}
wire w169;    //: /sn:0 {0}(1,1)(1,1){1}
wire w857;    //: /sn:0 {0}(1,1)(1,1){1}
wire w714;    //: /sn:0 {0}(1,1)(1,1){1}
wire w132;    //: /sn:0 {0}(1,1)(1,1){1}
wire w723;    //: /sn:0 {0}(1,1)(1,1){1}
wire w65;    //: /sn:0 {0}(1,1)(1,1){1}
wire w794;    //: /sn:0 {0}(1,1)(1,1){1}
wire w92;    //: /sn:0 {0}(1,1)(1,1){1}
wire w456;    //: /sn:0 {0}(1,1)(1,1){1}
wire w308;    //: /sn:0 {0}(1,1)(1,1){1}
wire w162;    //: /sn:0 {0}(1,1)(1,1){1}
wire w222;    //: /sn:0 {0}(1,1)(1,1){1}
wire w877;    //: /sn:0 {0}(1,1)(1,1){1}
wire w946;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1002;    //: /sn:0 {0}(1,1)(1,1){1}
wire w381;    //: /sn:0 {0}(1,1)(1,1){1}
wire w286;    //: /sn:0 {0}(1,1)(1,1){1}
wire w636;    //: /sn:0 {0}(1,1)(1,1){1}
wire w762;    //: /sn:0 {0}(1,1)(1,1){1}
wire w318;    //: /sn:0 {0}(1,1)(1,1){1}
wire w173;    //: /sn:0 {0}(1,1)(1,1){1}
wire w252;    //: /sn:0 {0}(1,1)(1,1){1}
wire w105;    //: /sn:0 {0}(1,1)(1,1){1}
wire w148;    //: /sn:0 {0}(1,1)(1,1){1}
wire w604;    //: /sn:0 {0}(1,1)(1,1){1}
wire w860;    //: /sn:0 {0}(1,1)(1,1){1}
wire w72;    //: /sn:0 {0}(1,1)(1,1){1}
wire w817;    //: /sn:0 {0}(1,1)(1,1){1}
wire w33;    //: /sn:0 {0}(1,1)(1,1){1}
wire w863;    //: /sn:0 {0}(1,1)(1,1){1}
wire w384;    //: /sn:0 {0}(1,1)(1,1){1}
wire w503;    //: /sn:0 {0}(1,1)(1,1){1}
wire w800;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1008;    //: /sn:0 {0}(1,1)(1,1){1}
wire w981;    //: /sn:0 {0}(1,1)(1,1){1}
wire w423;    //: /sn:0 {0}(1,1)(1,1){1}
wire w219;    //: /sn:0 {0}(1,1)(1,1){1}
wire w145;    //: /sn:0 {0}(1,1)(1,1){1}
wire w305;    //: /sn:0 {0}(1,1)(1,1){1}
wire w39;    //: /sn:0 {0}(1,1)(1,1){1}
wire w909;    //: /sn:0 {0}(1,1)(1,1){1}
wire w166;    //: /sn:0 {0}(1,1)(1,1){1}
wire w386;    //: /sn:0 {0}(1,1)(1,1){1}
wire w14;    //: /sn:0 {0}(1,1)(1,1){1}
wire w141;    //: /sn:0 {0}(1,1)(1,1){1}
wire w195;    //: /sn:0 {0}(1,1)(1,1){1}
wire w874;    //: /sn:0 {0}(1,1)(1,1){1}
wire w292;    //: /sn:0 {0}(1,1)(1,1){1}
wire w182;    //: /sn:0 {0}(1,1)(1,1){1}
wire w302;    //: /sn:0 {0}(1,1)(1,1){1}
wire w194;    //: /sn:0 {0}(1,1)(1,1){1}
wire w128;    //: /sn:0 {0}(1,1)(1,1){1}
wire w939;    //: /sn:0 {0}(1,1)(1,1){1}
wire w558;    //: /sn:0 {0}(1,1)(1,1){1}
wire w898;    //: /sn:0 {0}(1,1)(1,1){1}
wire w389;    //: /sn:0 {0}(1,1)(1,1){1}
wire w360;    //: /sn:0 {0}(1,1)(1,1){1}
wire w284;    //: /sn:0 {0}(1,1)(1,1){1}
wire w774;    //: /sn:0 {0}(1,1)(1,1){1}
wire w887;    //: /sn:0 {0}(1,1)(1,1){1}
wire w276;    //: /sn:0 {0}(1,1)(1,1){1}
wire w701;    //: /sn:0 {0}(1,1)(1,1){1}
wire w708;    //: /sn:0 {0}(1,1)(1,1){1}
wire w992;    //: /sn:0 {0}(1,1)(1,1){1}
wire w989;    //: /sn:0 {0}(1,1)(1,1){1}
wire w41;    //: /sn:0 {0}(1,1)(1,1){1}
wire w533;    //: /sn:0 {0}(1,1)(1,1){1}
wire w324;    //: /sn:0 {0}(1,1)(1,1){1}
wire w740;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1000;    //: /sn:0 {0}(1,1)(1,1){1}
wire w888;    //: /sn:0 {0}(1,1)(1,1){1}
wire w967;    //: /sn:0 {0}(1,1)(1,1){1}
wire w467;    //: /sn:0 {0}(1,1)(1,1){1}
wire w791;    //: /sn:0 {0}(1,1)(1,1){1}
wire w813;    //: /sn:0 {0}(1,1)(1,1){1}
wire w258;    //: /sn:0 {0}(1,1)(1,1){1}
wire w648;    //: /sn:0 {0}(1,1)(1,1){1}
wire w908;    //: /sn:0 {0}(1,1)(1,1){1}
wire w728;    //: /sn:0 {0}(1,1)(1,1){1}
wire w382;    //: /sn:0 {0}(1,1)(1,1){1}
wire w192;    //: /sn:0 {0}(1,1)(1,1){1}
wire w465;    //: /sn:0 {0}(1,1)(1,1){1}
wire w22;    //: /sn:0 {0}(1,1)(1,1){1}
wire w660;    //: /sn:0 {0}(1,1)(1,1){1}
wire w117;    //: /sn:0 {0}(1,1)(1,1){1}
wire w555;    //: /sn:0 {0}(1,1)(1,1){1}
wire w172;    //: /sn:0 {0}(1,1)(1,1){1}
wire w893;    //: /sn:0 {0}(1,1)(1,1){1}
wire w401;    //: /sn:0 {0}(1,1)(1,1){1}
wire w771;    //: /sn:0 {0}(1,1)(1,1){1}
wire w542;    //: /sn:0 {0}(1,1)(1,1){1}
wire w200;    //: /sn:0 {0}(1,1)(1,1){1}
wire w620;    //: /sn:0 {0}(1,1)(1,1){1}
wire w411;    //: /sn:0 {0}(1,1)(1,1){1}
wire w792;    //: /sn:0 {0}(1,1)(1,1){1}
wire w231;    //: /sn:0 {0}(1,1)(1,1){1}
wire w878;    //: /sn:0 {0}(1,1)(1,1){1}
wire w443;    //: /sn:0 {0}(1,1)(1,1){1}
wire w264;    //: /sn:0 {0}(1,1)(1,1){1}
wire w707;    //: /sn:0 {0}(1,1)(1,1){1}
wire w952;    //: /sn:0 {0}(1,1)(1,1){1}
wire w421;    //: /sn:0 {0}(1,1)(1,1){1}
wire w370;    //: /sn:0 {0}(1,1)(1,1){1}
wire w678;    //: /sn:0 {0}(1,1)(1,1){1}
wire w495;    //: /sn:0 {0}(1,1)(1,1){1}
wire w394;    //: /sn:0 {0}(1,1)(1,1){1}
wire w60;    //: /sn:0 {0}(1,1)(1,1){1}
wire w486;    //: /sn:0 {0}(1,1)(1,1){1}
wire w790;    //: /sn:0 {0}(1,1)(1,1){1}
wire w996;    //: /sn:0 {0}(1,1)(1,1){1}
wire w931;    //: /sn:0 {0}(1,1)(1,1){1}
wire w15;    //: /sn:0 {0}(1,1)(1,1){1}
wire w494;    //: /sn:0 {0}(1,1)(1,1){1}
wire w731;    //: /sn:0 {0}(1,1)(1,1){1}
wire w535;    //: /sn:0 {0}(1,1)(1,1){1}
wire w560;    //: /sn:0 {0}(1,1)(1,1){1}
wire w634;    //: /sn:0 {0}(1,1)(1,1){1}
wire w109;    //: /sn:0 {0}(1,1)(1,1){1}
wire w567;    //: /sn:0 {0}(1,1)(1,1){1}
wire w615;    //: /sn:0 {0}(1,1)(1,1){1}
wire w619;    //: /sn:0 {0}(1,1)(1,1){1}
wire w979;    //: /sn:0 {0}(1,1)(1,1){1}
wire w97;    //: /sn:0 {0}(1,1)(1,1){1}
wire w114;    //: /sn:0 {0}(1,1)(1,1){1}
wire w261;    //: /sn:0 {0}(1,1)(1,1){1}
wire w245;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1010;    //: /sn:0 {0}(1,1)(1,1){1}
wire w480;    //: /sn:0 {0}(1,1)(1,1){1}
wire w705;    //: /sn:0 {0}(1,1)(1,1){1}
wire w836;    //: /sn:0 {0}(1,1)(1,1){1}
wire w617;    //: /sn:0 {0}(1,1)(1,1){1}
wire w940;    //: /sn:0 {0}(1,1)(1,1){1}
wire w957;    //: /sn:0 {0}(1,1)(1,1){1}
wire w521;    //: /sn:0 {0}(1,1)(1,1){1}
wire w391;    //: /sn:0 {0}(1,1)(1,1){1}
wire w24;    //: /sn:0 {0}(1,1)(1,1){1}
wire w221;    //: /sn:0 {0}(1,1)(1,1){1}
wire w140;    //: /sn:0 {0}(1,1)(1,1){1}
wire w822;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1022;    //: /sn:0 {0}(1,1)(1,1){1}
wire w372;    //: /sn:0 {0}(1,1)(1,1){1}
wire w227;    //: /sn:0 {0}(1,1)(1,1){1}
wire w243;    //: /sn:0 {0}(1,1)(1,1){1}
wire w212;    //: /sn:0 {0}(1,1)(1,1){1}
wire w18;    //: /sn:0 {0}(1,1)(1,1){1}
wire w118;    //: /sn:0 {0}(1,1)(1,1){1}
wire w722;    //: /sn:0 {0}(1,1)(1,1){1}
wire w808;    //: /sn:0 {0}(1,1)(1,1){1}
wire w865;    //: /sn:0 {0}(1,1)(1,1){1}
wire w363;    //: /sn:0 {0}(1,1)(1,1){1}
wire w164;    //: /sn:0 {0}(1,1)(1,1){1}
wire w464;    //: /sn:0 {0}(1,1)(1,1){1}
wire w732;    //: /sn:0 {0}(1,1)(1,1){1}
wire w407;    //: /sn:0 {0}(1,1)(1,1){1}
wire w451;    //: /sn:0 {0}(1,1)(1,1){1}
wire w595;    //: /sn:0 {0}(1,1)(1,1){1}
wire w639;    //: /sn:0 {0}(1,1)(1,1){1}
wire w59;    //: /sn:0 {0}(1,1)(1,1){1}
wire w525;    //: /sn:0 {0}(1,1)(1,1){1}
wire w62;    //: /sn:0 {0}(1,1)(1,1){1}
wire w588;    //: /sn:0 {0}(1,1)(1,1){1}
wire w602;    //: /sn:0 {0}(1,1)(1,1){1}
wire w624;    //: /sn:0 {0}(1,1)(1,1){1}
wire w787;    //: /sn:0 {0}(1,1)(1,1){1}
wire w853;    //: /sn:0 {0}(1,1)(1,1){1}
wire w150;    //: /sn:0 {0}(1,1)(1,1){1}
wire w189;    //: /sn:0 {0}(1,1)(1,1){1}
wire w206;    //: /sn:0 {0}(1,1)(1,1){1}
wire w353;    //: /sn:0 {0}(1,1)(1,1){1}
wire w354;    //: /sn:0 {0}(1,1)(1,1){1}
wire w918;    //: /sn:0 {0}(1,1)(1,1){1}
wire w325;    //: /sn:0 {0}(1,1)(1,1){1}
wire w569;    //: /sn:0 {0}(1,1)(1,1){1}
wire w809;    //: /sn:0 {0}(1,1)(1,1){1}
wire w796;    //: /sn:0 {0}(1,1)(1,1){1}
wire w945;    //: /sn:0 {0}(1,1)(1,1){1}
wire w879;    //: /sn:0 {0}(1,1)(1,1){1}
wire w784;    //: /sn:0 {0}(1,1)(1,1){1}
wire w404;    //: /sn:0 {0}(1,1)(1,1){1}
wire w218;    //: /sn:0 {0}(1,1)(1,1){1}
wire w56;    //: /sn:0 {0}(1,1)(1,1){1}
wire w804;    //: /sn:0 {0}(1,1)(1,1){1}
wire w876;    //: /sn:0 {0}(1,1)(1,1){1}
wire w962;    //: /sn:0 {0}(1,1)(1,1){1}
wire w376;    //: /sn:0 {0}(1,1)(1,1){1}
wire w183;    //: /sn:0 {0}(1,1)(1,1){1}
wire w628;    //: /sn:0 {0}(1,1)(1,1){1}
wire w663;    //: /sn:0 {0}(1,1)(1,1){1}
wire w383;    //: /sn:0 {0}(1,1)(1,1){1}
wire w120;    //: /sn:0 {0}(1,1)(1,1){1}
wire w572;    //: /sn:0 {0}(1,1)(1,1){1}
wire w676;    //: /sn:0 {0}(1,1)(1,1){1}
wire w677;    //: /sn:0 {0}(1,1)(1,1){1}
wire w168;    //: /sn:0 {0}(1,1)(1,1){1}
wire w849;    //: /sn:0 {0}(1,1)(1,1){1}
wire w327;    //: /sn:0 {0}(1,1)(1,1){1}
wire w54;    //: /sn:0 {0}(1,1)(1,1){1}
wire w399;    //: /sn:0 {0}(1,1)(1,1){1}
wire w632;    //: /sn:0 {0}(1,1)(1,1){1}
wire w734;    //: /sn:0 {0}(1,1)(1,1){1}
wire w445;    //: /sn:0 {0}(1,1)(1,1){1}
wire w20;    //: /sn:0 {0}(1,1)(1,1){1}
wire w124;    //: /sn:0 {0}(1,1)(1,1){1}
wire w606;    //: /sn:0 {0}(1,1)(1,1){1}
wire w687;    //: /sn:0 {0}(1,1)(1,1){1}
wire w950;    //: /sn:0 {0}(1,1)(1,1){1}
wire w763;    //: /sn:0 {0}(1,1)(1,1){1}
wire w507;    //: /sn:0 {0}(1,1)(1,1){1}
wire w437;    //: /sn:0 {0}(1,1)(1,1){1}
wire w125;    //: /sn:0 {0}(1,1)(1,1){1}
wire w929;    //: /sn:0 {0}(1,1)(1,1){1}
wire w393;    //: /sn:0 {0}(1,1)(1,1){1}
wire w17;    //: /sn:0 {0}(1,1)(1,1){1}
wire w599;    //: /sn:0 {0}(1,1)(1,1){1}
wire w53;    //: /sn:0 {0}(1,1)(1,1){1}
wire w263;    //: /sn:0 {0}(1,1)(1,1){1}
wire w633;    //: /sn:0 {0}(1,1)(1,1){1}
wire w649;    //: /sn:0 {0}(1,1)(1,1){1}
wire w113;    //: /sn:0 {0}(1,1)(1,1){1}
wire w515;    //: /sn:0 {0}(1,1)(1,1){1}
wire w262;    //: /sn:0 {0}(1,1)(1,1){1}
wire w224;    //: /sn:0 {0}(1,1)(1,1){1}
wire w273;    //: /sn:0 {0}(1,1)(1,1){1}
wire w438;    //: /sn:0 {0}(1,1)(1,1){1}
wire w388;    //: /sn:0 {0}(1,1)(1,1){1}
wire w188;    //: /sn:0 {0}(1,1)(1,1){1}
wire w187;    //: /sn:0 {0}(1,1)(1,1){1}
wire w783;    //: /sn:0 {0}(1,1)(1,1){1}
wire w548;    //: /sn:0 {0}(1,1)(1,1){1}
wire w735;    //: /sn:0 {0}(1,1)(1,1){1}
wire w773;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1009;    //: /sn:0 {0}(1,1)(1,1){1}
wire w432;    //: /sn:0 {0}(1,1)(1,1){1}
wire w6;    //: /sn:0 {0}(1,1)(1,1){1}
wire w7;    //: /sn:0 {0}(1,1)(1,1){1}
wire w61;    //: /sn:0 {0}(1,1)(1,1){1}
wire w99;    //: /sn:0 {0}(1,1)(1,1){1}
wire w609;    //: /sn:0 {0}(1,1)(1,1){1}
wire w751;    //: /sn:0 {0}(1,1)(1,1){1}
wire w380;    //: /sn:0 {0}(1,1)(1,1){1}
wire w352;    //: /sn:0 {0}(1,1)(1,1){1}
wire w531;    //: /sn:0 {0}(1,1)(1,1){1}
wire w349;    //: /sn:0 {0}(1,1)(1,1){1}
wire w106;    //: /sn:0 {0}(1,1)(1,1){1}
wire w652;    //: /sn:0 {0}(1,1)(1,1){1}
wire w718;    //: /sn:0 {0}(1,1)(1,1){1}
wire w743;    //: /sn:0 {0}(1,1)(1,1){1}
wire w984;    //: /sn:0 {0}(1,1)(1,1){1}
wire w356;    //: /sn:0 {0}(1,1)(1,1){1}
wire w43;    //: /sn:0 {0}(1,1)(1,1){1}
wire w476;    //: /sn:0 {0}(1,1)(1,1){1}
wire w672;    //: /sn:0 {0}(1,1)(1,1){1}
wire w847;    //: /sn:0 {0}(1,1)(1,1){1}
wire w907;    //: /sn:0 {0}(1,1)(1,1){1}
wire w58;    //: /sn:0 {0}(1,1)(1,1){1}
wire w697;    //: /sn:0 {0}(1,1)(1,1){1}
wire w772;    //: /sn:0 {0}(1,1)(1,1){1}
wire w781;    //: /sn:0 {0}(1,1)(1,1){1}
wire w629;    //: /sn:0 {0}(1,1)(1,1){1}
wire w844;    //: /sn:0 {0}(1,1)(1,1){1}
wire w971;    //: /sn:0 {0}(1,1)(1,1){1}
wire w184;    //: /sn:0 {0}(1,1)(1,1){1}
wire w662;    //: /sn:0 {0}(1,1)(1,1){1}
wire w283;    //: /sn:0 {0}(1,1)(1,1){1}
wire w830;    //: /sn:0 {0}(1,1)(1,1){1}
wire w958;    //: /sn:0 {0}(1,1)(1,1){1}
wire w703;    //: /sn:0 {0}(1,1)(1,1){1}
wire w758;    //: /sn:0 {0}(1,1)(1,1){1}
wire w834;    //: /sn:0 {0}(1,1)(1,1){1}
wire w165;    //: /sn:0 {0}(1,1)(1,1){1}
wire w713;    //: /sn:0 {0}(1,1)(1,1){1}
wire w819;    //: /sn:0 {0}(1,1)(1,1){1}
wire w57;    //: /sn:0 {0}(1,1)(1,1){1}
wire w136;    //: /sn:0 {0}(1,1)(1,1){1}
wire w910;    //: /sn:0 {0}(1,1)(1,1){1}
wire w610;    //: /sn:0 {0}(1,1)(1,1){1}
wire w505;    //: /sn:0 {0}(1,1)(1,1){1}
wire w94;    //: /sn:0 {0}(1,1)(1,1){1}
wire w561;    //: /sn:0 {0}(1,1)(1,1){1}
wire w754;    //: /sn:0 {0}(1,1)(1,1){1}
wire w960;    //: /sn:0 {0}(1,1)(1,1){1}
wire w440;    //: /sn:0 {0}(1,1)(1,1){1}
wire w904;    //: /sn:0 {0}(1,1)(1,1){1}
wire w337;    //: /sn:0 {0}(1,1)(1,1){1}
wire w201;    //: /sn:0 {0}(1,1)(1,1){1}
wire w685;    //: /sn:0 {0}(1,1)(1,1){1}
wire w727;    //: /sn:0 {0}(1,1)(1,1){1}
wire w459;    //: /sn:0 {0}(1,1)(1,1){1}
wire w553;    //: /sn:0 {0}(1,1)(1,1){1}
wire w613;    //: /sn:0 {0}(1,1)(1,1){1}
wire w122;    //: /sn:0 {0}(1,1)(1,1){1}
wire w826;    //: /sn:0 {0}(1,1)(1,1){1}
wire w944;    //: /sn:0 {0}(1,1)(1,1){1}
wire w220;    //: /sn:0 {0}(1,1)(1,1){1}
wire w250;    //: /sn:0 {0}(1,1)(1,1){1}
wire w38;    //: /sn:0 {0}(1,1)(1,1){1}
wire w845;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1013;    //: /sn:0 {0}(1,1)(1,1){1}
wire w977;    //: /sn:0 {0}(1,1)(1,1){1}
wire w3;    //: /sn:0 {0}(1,1)(1,1){1}
wire w408;    //: /sn:0 {0}(1,1)(1,1){1}
wire w127;    //: /sn:0 {0}(1,1)(1,1){1}
wire w493;    //: /sn:0 {0}(1,1)(1,1){1}
wire w133;    //: /sn:0 {0}(1,1)(1,1){1}
wire w635;    //: /sn:0 {0}(1,1)(1,1){1}
wire w75;    //: /sn:0 {0}(1,1)(1,1){1}
wire w757;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1006;    //: /sn:0 {0}(1,1)(1,1){1}
wire w209;    //: /sn:0 {0}(1,1)(1,1){1}
wire w502;    //: /sn:0 {0}(1,1)(1,1){1}
wire w564;    //: /sn:0 {0}(1,1)(1,1){1}
wire w420;    //: /sn:0 {0}(1,1)(1,1){1}
wire w215;    //: /sn:0 {0}(1,1)(1,1){1}
wire w529;    //: /sn:0 {0}(1,1)(1,1){1}
wire w706;    //: /sn:0 {0}(1,1)(1,1){1}
wire w975;    //: /sn:0 {0}(1,1)(1,1){1}
wire w36;    //: /sn:0 {0}(1,1)(1,1){1}
wire w496;    //: /sn:0 {0}(1,1)(1,1){1}
wire w472;    //: /sn:0 {0}(1,1)(1,1){1}
wire w419;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1019;    //: /sn:0 {0}(1,1)(1,1){1}
wire w82;    //: /sn:0 {0}(1,1)(1,1){1}
wire w303;    //: /sn:0 {0}(1,1)(1,1){1}
wire w158;    //: /sn:0 {0}(1,1)(1,1){1}
wire w650;    //: /sn:0 {0}(1,1)(1,1){1}
wire w571;    //: /sn:0 {0}(1,1)(1,1){1}
wire w439;    //: /sn:0 {0}(1,1)(1,1){1}
wire w711;    //: /sn:0 {0}(1,1)(1,1){1}
wire w748;    //: /sn:0 {0}(1,1)(1,1){1}
wire w296;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1017;    //: /sn:0 {0}(1,1)(1,1){1}
wire w449;    //: /sn:0 {0}(1,1)(1,1){1}
wire w402;    //: /sn:0 {0}(1,1)(1,1){1}
wire w802;    //: /sn:0 {0}(1,1)(1,1){1}
wire w749;    //: /sn:0 {0}(1,1)(1,1){1}
wire w875;    //: /sn:0 {0}(1,1)(1,1){1}
wire w978;    //: /sn:0 {0}(1,1)(1,1){1}
wire w398;    //: /sn:0 {0}(1,1)(1,1){1}
wire w226;    //: /sn:0 {0}(1,1)(1,1){1}
wire w301;    //: /sn:0 {0}(1,1)(1,1){1}
wire w78;    //: /sn:0 {0}(1,1)(1,1){1}
wire w479;    //: /sn:0 {0}(1,1)(1,1){1}
wire w517;    //: /sn:0 {0}(1,1)(1,1){1}
wire w608;    //: /sn:0 {0}(1,1)(1,1){1}
wire w715;    //: /sn:0 {0}(1,1)(1,1){1}
wire w998;    //: /sn:0 {0}(1,1)(1,1){1}
wire w246;    //: /sn:0 {0}(1,1)(1,1){1}
wire w86;    //: /sn:0 {0}(1,1)(1,1){1}
wire w138;    //: /sn:0 {0}(1,1)(1,1){1}
wire w544;    //: /sn:0 {0}(1,1)(1,1){1}
wire w29;    //: /sn:0 {0}(1,1)(1,1){1}
wire w80;    //: /sn:0 {0}(1,1)(1,1){1}
wire w949;    //: /sn:0 {0}(1,1)(1,1){1}
wire w42;    //: /sn:0 {0}(1,1)(1,1){1}
wire w147;    //: /sn:0 {0}(1,1)(1,1){1}
wire w793;    //: /sn:0 {0}(1,1)(1,1){1}
wire w825;    //: /sn:0 {0}(1,1)(1,1){1}
wire w317;    //: /sn:0 {0}(1,1)(1,1){1}
wire w892;    //: /sn:0 {0}(1,1)(1,1){1}
wire w976;    //: /sn:0 {0}(1,1)(1,1){1}
wire w46;    //: /sn:0 {0}(1,1)(1,1){1}
wire w175;    //: /sn:0 {0}(1,1)(1,1){1}
wire w530;    //: /sn:0 {0}(1,1)(1,1){1}
wire w645;    //: /sn:0 {0}(1,1)(1,1){1}
wire w721;    //: /sn:0 {0}(1,1)(1,1){1}
wire w885;    //: /sn:0 {0}(1,1)(1,1){1}
wire w578;    //: /sn:0 {0}(1,1)(1,1){1}
wire w959;    //: /sn:0 {0}(1,1)(1,1){1}
wire w291;    //: /sn:0 {0}(1,1)(1,1){1}
wire w638;    //: /sn:0 {0}(1,1)(1,1){1}
wire w871;    //: /sn:0 {0}(1,1)(1,1){1}
wire w675;    //: /sn:0 {0}(1,1)(1,1){1}
wire w937;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1007;    //: /sn:0 {0}(1,1)(1,1){1}
wire w229;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1001;    //: /sn:0 {0}(1,1)(1,1){1}
wire w285;    //: /sn:0 {0}(1,1)(1,1){1}
wire w64;    //: /sn:0 {0}(1,1)(1,1){1}
wire w868;    //: /sn:0 {0}(1,1)(1,1){1}
wire w575;    //: /sn:0 {0}(1,1)(1,1){1}
wire w644;    //: /sn:0 {0}(1,1)(1,1){1}
wire w756;    //: /sn:0 {0}(1,1)(1,1){1}
wire w374;    //: /sn:0 {0}(1,1)(1,1){1}
wire w988;    //: /sn:0 {0}(1,1)(1,1){1}
wire w603;    //: /sn:0 {0}(1,1)(1,1){1}
wire w693;    //: /sn:0 {0}(1,1)(1,1){1}
wire w31;    //: /sn:0 {0}(1,1)(1,1){1}
wire w100;    //: /sn:0 {0}(1,1)(1,1){1}
wire w251;    //: /sn:0 {0}(1,1)(1,1){1}
wire w161;    //: /sn:0 {0}(1,1)(1,1){1}
wire w991;    //: /sn:0 {0}(1,1)(1,1){1}
wire w334;    //: /sn:0 {0}(1,1)(1,1){1}
wire w235;    //: /sn:0 {0}(1,1)(1,1){1}
wire w196;    //: /sn:0 {0}(1,1)(1,1){1}
wire w346;    //: /sn:0 {0}(1,1)(1,1){1}
wire w205;    //: /sn:0 {0}(1,1)(1,1){1}
wire w154;    //: /sn:0 {0}(1,1)(1,1){1}
wire w782;    //: /sn:0 {0}(1,1)(1,1){1}
wire w815;    //: /sn:0 {0}(1,1)(1,1){1}
wire w953;    //: /sn:0 {0}(1,1)(1,1){1}
wire w466;    //: /sn:0 {0}(1,1)(1,1){1}
wire w422;    //: /sn:0 {0}(1,1)(1,1){1}
wire w68;    //: /sn:0 {0}(1,1)(1,1){1}
wire w938;    //: /sn:0 {0}(1,1)(1,1){1}
wire w867;    //: /sn:0 {0}(1,1)(1,1){1}
wire w85;    //: /sn:0 {0}(1,1)(1,1){1}
wire w197;    //: /sn:0 {0}(1,1)(1,1){1}
wire w110;    //: /sn:0 {0}(1,1)(1,1){1}
wire w651;    //: /sn:0 {0}(1,1)(1,1){1}
wire w785;    //: /sn:0 {0}(1,1)(1,1){1}
wire w446;    //: /sn:0 {0}(1,1)(1,1){1}
wire w48;    //: /sn:0 {0}(1,1)(1,1){1}
wire w5;    //: /sn:0 {0}(1,1)(1,1){1}
wire w667;    //: /sn:0 {0}(1,1)(1,1){1}
wire w828;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1015;    //: /sn:0 {0}(1,1)(1,1){1}
wire w342;    //: /sn:0 {0}(1,1)(1,1){1}
wire w26;    //: /sn:0 {0}(1,1)(1,1){1}
wire w630;    //: /sn:0 {0}(1,1)(1,1){1}
wire w364;    //: /sn:0 {0}(1,1)(1,1){1}
wire w270;    //: /sn:0 {0}(1,1)(1,1){1}
wire w780;    //: /sn:0 {0}(1,1)(1,1){1}
wire w73;    //: /sn:0 {0}(1,1)(1,1){1}
wire w96;    //: /sn:0 {0}(1,1)(1,1){1}
wire w955;    //: /sn:0 {0}(1,1)(1,1){1}
wire w405;    //: /sn:0 {0}(1,1)(1,1){1}
wire w359;    //: /sn:0 {0}(1,1)(1,1){1}
wire w339;    //: /sn:0 {0}(1,1)(1,1){1}
wire w320;    //: /sn:0 {0}(1,1)(1,1){1}
wire w244;    //: /sn:0 {0}(1,1)(1,1){1}
wire w16;    //: /sn:0 {0}(1,1)(1,1){1}
wire w963;    //: /sn:0 {0}(1,1)(1,1){1}
wire w387;    //: /sn:0 {0}(1,1)(1,1){1}
wire w81;    //: /sn:0 {0}(1,1)(1,1){1}
wire w89;    //: /sn:0 {0}(1,1)(1,1){1}
wire w576;    //: /sn:0 {0}(1,1)(1,1){1}
wire w616;    //: /sn:0 {0}(1,1)(1,1){1}
wire w518;    //: /sn:0 {0}(1,1)(1,1){1}
wire w689;    //: /sn:0 {0}(1,1)(1,1){1}
wire w899;    //: /sn:0 {0}(1,1)(1,1){1}
wire w417;    //: /sn:0 {0}(1,1)(1,1){1}
wire w0;    //: /sn:0 {0}(1,1)(1,1){1}
wire w313;    //: /sn:0 {0}(1,1)(1,1){1}
wire w240;    //: /sn:0 {0}(1,1)(1,1){1}
wire w233;    //: /sn:0 {0}(1,1)(1,1){1}
wire w987;    //: /sn:0 {0}(1,1)(1,1){1}
wire w926;    //: /sn:0 {0}(1,1)(1,1){1}
wire w287;    //: /sn:0 {0}(1,1)(1,1){1}
wire w956;    //: /sn:0 {0}(1,1)(1,1){1}
wire w934;    //: /sn:0 {0}(1,1)(1,1){1}
wire w176;    //: /sn:0 {0}(1,1)(1,1){1}
wire w691;    //: /sn:0 {0}(1,1)(1,1){1}
wire w745;    //: /sn:0 {0}(1,1)(1,1){1}
wire w866;    //: /sn:0 {0}(1,1)(1,1){1}
wire w919;    //: /sn:0 {0}(1,1)(1,1){1}
wire w770;    //: /sn:0 {0}(1,1)(1,1){1}
wire w23;    //: /sn:0 {0}(1,1)(1,1){1}
wire w174;    //: /sn:0 {0}(1,1)(1,1){1}
wire w671;    //: /sn:0 {0}(1,1)(1,1){1}
wire w859;    //: /sn:0 {0}(1,1)(1,1){1}
wire w225;    //: /sn:0 {0}(1,1)(1,1){1}
wire w506;    //: /sn:0 {0}(1,1)(1,1){1}
wire w556;    //: /sn:0 {0}(1,1)(1,1){1}
wire w811;    //: /sn:0 {0}(1,1)(1,1){1}
wire w547;    //: /sn:0 {0}(1,1)(1,1){1}
wire w589;    //: /sn:0 {0}(1,1)(1,1){1}
wire w725;    //: /sn:0 {0}(1,1)(1,1){1}
wire w71;    //: /sn:0 {0}(1,1)(1,1){1}
wire w559;    //: /sn:0 {0}(1,1)(1,1){1}
wire w948;    //: /sn:0 {0}(1,1)(1,1){1}
wire w400;    //: /sn:0 {0}(1,1)(1,1){1}
wire w492;    //: /sn:0 {0}(1,1)(1,1){1}
wire w851;    //: /sn:0 {0}(1,1)(1,1){1}
wire w255;    //: /sn:0 {0}(1,1)(1,1){1}
wire w710;    //: /sn:0 {0}(1,1)(1,1){1}
wire w742;    //: /sn:0 {0}(1,1)(1,1){1}
wire w900;    //: /sn:0 {0}(1,1)(1,1){1}
wire w345;    //: /sn:0 {0}(1,1)(1,1){1}
wire w2;    //: /sn:0 {0}(1,1)(1,1){1}
wire w77;    //: /sn:0 {0}(1,1)(1,1){1}
wire w570;    //: /sn:0 {0}(1,1)(1,1){1}
wire w366;    //: /sn:0 {0}(1,1)(1,1){1}
wire w601;    //: /sn:0 {0}(1,1)(1,1){1}
wire w943;    //: /sn:0 {0}(1,1)(1,1){1}
wire w289;    //: /sn:0 {0}(1,1)(1,1){1}
wire w190;    //: /sn:0 {0}(1,1)(1,1){1}
wire w778;    //: /sn:0 {0}(1,1)(1,1){1}
wire w897;    //: /sn:0 {0}(1,1)(1,1){1}
wire w562;    //: /sn:0 {0}(1,1)(1,1){1}
wire w679;    //: /sn:0 {0}(1,1)(1,1){1}
wire w839;    //: /sn:0 {0}(1,1)(1,1){1}
wire w142;    //: /sn:0 {0}(1,1)(1,1){1}
wire w155;    //: /sn:0 {0}(1,1)(1,1){1}
wire w509;    //: /sn:0 {0}(1,1)(1,1){1}
wire w50;    //: /sn:0 {0}(1,1)(1,1){1}
wire w970;    //: /sn:0 {0}(1,1)(1,1){1}
wire w527;    //: /sn:0 {0}(1,1)(1,1){1}
wire w453;    //: /sn:0 {0}(1,1)(1,1){1}
wire w927;    //: /sn:0 {0}(1,1)(1,1){1}
wire w93;    //: /sn:0 {0}(1,1)(1,1){1}
wire w816;    //: /sn:0 {0}(1,1)(1,1){1}
wire w983;    //: /sn:0 {0}(1,1)(1,1){1}
wire w135;    //: /sn:0 {0}(1,1)(1,1){1}
wire w625;    //: /sn:0 {0}(1,1)(1,1){1}
wire w216;    //: /sn:0 {0}(1,1)(1,1){1}
wire w425;    //: /sn:0 {0}(1,1)(1,1){1}
wire w288;    //: /sn:0 {0}(1,1)(1,1){1}
wire w753;    //: /sn:0 {0}(1,1)(1,1){1}
wire w429;    //: /sn:0 {0}(1,1)(1,1){1}
wire w373;    //: /sn:0 {0}(1,1)(1,1){1}
wire w750;    //: /sn:0 {0}(1,1)(1,1){1}
wire w357;    //: /sn:0 {0}(1,1)(1,1){1}
wire w37;    //: /sn:0 {0}(1,1)(1,1){1}
wire w843;    //: /sn:0 {0}(1,1)(1,1){1}
wire w34;    //: /sn:0 {0}(1,1)(1,1){1}
wire w688;    //: /sn:0 {0}(1,1)(1,1){1}
wire w820;    //: /sn:0 {0}(1,1)(1,1){1}
wire w254;    //: /sn:0 {0}(1,1)(1,1){1}
wire w102;    //: /sn:0 {0}(1,1)(1,1){1}
wire w157;    //: /sn:0 {0}(1,1)(1,1){1}
wire w593;    //: /sn:0 {0}(1,1)(1,1){1}
wire w475;    //: /sn:0 {0}(1,1)(1,1){1}
wire w917;    //: /sn:0 {0}(1,1)(1,1){1}
wire w673;    //: /sn:0 {0}(1,1)(1,1){1}
wire w724;    //: /sn:0 {0}(1,1)(1,1){1}
wire w435;    //: /sn:0 {0}(1,1)(1,1){1}
wire w886;    //: /sn:0 {0}(1,1)(1,1){1}
wire w668;    //: /sn:0 {0}(1,1)(1,1){1}
wire w269;    //: /sn:0 {0}(1,1)(1,1){1}
wire w511;    //: /sn:0 {0}(1,1)(1,1){1}
wire w210;    //: /sn:0 {0}(1,1)(1,1){1}
wire w747;    //: /sn:0 {0}(1,1)(1,1){1}
wire w40;    //: /sn:0 {0}(1,1)(1,1){1}
wire w217;    //: /sn:0 {0}(1,1)(1,1){1}
wire w30;    //: /sn:0 {0}(1,1)(1,1){1}
wire w605;    //: /sn:0 {0}(1,1)(1,1){1}
wire w812;    //: /sn:0 {0}(1,1)(1,1){1}
wire w873;    //: /sn:0 {0}(1,1)(1,1){1}
wire w928;    //: /sn:0 {0}(1,1)(1,1){1}
wire w146;    //: /sn:0 {0}(1,1)(1,1){1}
wire w149;    //: /sn:0 {0}(1,1)(1,1){1}
wire w858;    //: /sn:0 {0}(1,1)(1,1){1}
wire w942;    //: /sn:0 {0}(1,1)(1,1){1}
wire w500;    //: /sn:0 {0}(1,1)(1,1){1}
wire w457;    //: /sn:0 {0}(1,1)(1,1){1}
wire w350;    //: /sn:0 {0}(1,1)(1,1){1}
wire w895;    //: /sn:0 {0}(1,1)(1,1){1}
wire w186;    //: /sn:0 {0}(1,1)(1,1){1}
wire w752;    //: /sn:0 {0}(1,1)(1,1){1}
wire w954;    //: /sn:0 {0}(1,1)(1,1){1}
wire w450;    //: /sn:0 {0}(1,1)(1,1){1}
wire w670;    //: /sn:0 {0}(1,1)(1,1){1}
wire w775;    //: /sn:0 {0}(1,1)(1,1){1}
wire w143;    //: /sn:0 {0}(1,1)(1,1){1}
wire w482;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1004;    //: /sn:0 {0}(1,1)(1,1){1}
wire w348;    //: /sn:0 {0}(1,1)(1,1){1}
wire w9;    //: /sn:0 {0}(1,1)(1,1){1}
wire w79;    //: /sn:0 {0}(1,1)(1,1){1}
wire w55;    //: /sn:0 {0}(1,1)(1,1){1}
wire w490;    //: /sn:0 {0}(1,1)(1,1){1}
wire w626;    //: /sn:0 {0}(1,1)(1,1){1}
wire w803;    //: /sn:0 {0}(1,1)(1,1){1}
wire w214;    //: /sn:0 {0}(1,1)(1,1){1}
wire w203;    //: /sn:0 {0}(1,1)(1,1){1}
wire w546;    //: /sn:0 {0}(1,1)(1,1){1}
wire w666;    //: /sn:0 {0}(1,1)(1,1){1}
wire w789;    //: /sn:0 {0}(1,1)(1,1){1}
wire w855;    //: /sn:0 {0}(1,1)(1,1){1}
wire w643;    //: /sn:0 {0}(1,1)(1,1){1}
wire w514;    //: /sn:0 {0}(1,1)(1,1){1}
wire w426;    //: /sn:0 {0}(1,1)(1,1){1}
wire w152;    //: /sn:0 {0}(1,1)(1,1){1}
wire w180;    //: /sn:0 {0}(1,1)(1,1){1}
wire w661;    //: /sn:0 {0}(1,1)(1,1){1}
wire w181;    //: /sn:0 {0}(1,1)(1,1){1}
wire w777;    //: /sn:0 {0}(1,1)(1,1){1}
wire w623;    //: /sn:0 {0}(1,1)(1,1){1}
wire w746;    //: /sn:0 {0}(1,1)(1,1){1}
wire w447;    //: /sn:0 {0}(1,1)(1,1){1}
wire w442;    //: /sn:0 {0}(1,1)(1,1){1}
wire w379;    //: /sn:0 {0}(1,1)(1,1){1}
wire w586;    //: /sn:0 {0}(1,1)(1,1){1}
wire w896;    //: /sn:0 {0}(1,1)(1,1){1}
wire w901;    //: /sn:0 {0}(1,1)(1,1){1}
wire w730;    //: /sn:0 {0}(1,1)(1,1){1}
wire w932;    //: /sn:0 {0}(1,1)(1,1){1}
wire w577;    //: /sn:0 {0}(1,1)(1,1){1}
wire w631;    //: /sn:0 {0}(1,1)(1,1){1}
wire w726;    //: /sn:0 {0}(1,1)(1,1){1}
wire w444;    //: /sn:0 {0}(1,1)(1,1){1}
wire w484;    //: /sn:0 {0}(1,1)(1,1){1}
wire w694;    //: /sn:0 {0}(1,1)(1,1){1}
wire w74;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1005;    //: /sn:0 {0}(1,1)(1,1){1}
wire w598;    //: /sn:0 {0}(1,1)(1,1){1}
wire w101;    //: /sn:0 {0}(1,1)(1,1){1}
wire w612;    //: /sn:0 {0}(1,1)(1,1){1}
wire w265;    //: /sn:0 {0}(1,1)(1,1){1}
wire w654;    //: /sn:0 {0}(1,1)(1,1){1}
wire w741;    //: /sn:0 {0}(1,1)(1,1){1}
wire w972;    //: /sn:0 {0}(1,1)(1,1){1}
wire w768;    //: /sn:0 {0}(1,1)(1,1){1}
wire w801;    //: /sn:0 {0}(1,1)(1,1){1}
wire w824;    //: /sn:0 {0}(1,1)(1,1){1}
wire w282;    //: /sn:0 {0}(1,1)(1,1){1}
wire w454;    //: /sn:0 {0}(1,1)(1,1){1}
wire w665;    //: /sn:0 {0}(1,1)(1,1){1}
wire w720;    //: /sn:0 {0}(1,1)(1,1){1}
wire w519;    //: /sn:0 {0}(1,1)(1,1){1}
wire w854;    //: /sn:0 {0}(1,1)(1,1){1}
wire w485;    //: /sn:0 {0}(1,1)(1,1){1}
wire w460;    //: /sn:0 {0}(1,1)(1,1){1}
wire w395;    //: /sn:0 {0}(1,1)(1,1){1}
wire w664;    //: /sn:0 {0}(1,1)(1,1){1}
wire w799;    //: /sn:0 {0}(1,1)(1,1){1}
wire w322;    //: /sn:0 {0}(1,1)(1,1){1}
wire w312;    //: /sn:0 {0}(1,1)(1,1){1}
wire w795;    //: /sn:0 {0}(1,1)(1,1){1}
wire w277;    //: /sn:0 {0}(1,1)(1,1){1}
wire w579;    //: /sn:0 {0}(1,1)(1,1){1}
wire w935;    //: /sn:0 {0}(1,1)(1,1){1}
wire w999;    //: /sn:0 {0}(1,1)(1,1){1}
wire w982;    //: /sn:0 {0}(1,1)(1,1){1}
wire w247;    //: /sn:0 {0}(1,1)(1,1){1}
wire w585;    //: /sn:0 {0}(1,1)(1,1){1}
wire w592;    //: /sn:0 {0}(1,1)(1,1){1}
wire w690;    //: /sn:0 {0}(1,1)(1,1){1}
wire w905;    //: /sn:0 {0}(1,1)(1,1){1}
wire w336;    //: /sn:0 {0}(1,1)(1,1){1}
wire w112;    //: /sn:0 {0}(1,1)(1,1){1}
wire w646;    //: /sn:0 {0}(1,1)(1,1){1}
wire w700;    //: /sn:0 {0}(1,1)(1,1){1}
wire w986;    //: /sn:0 {0}(1,1)(1,1){1}
wire w618;    //: /sn:0 {0}(1,1)(1,1){1}
wire w764;    //: /sn:0 {0}(1,1)(1,1){1}
wire w653;    //: /sn:0 {0}(1,1)(1,1){1}
wire w882;    //: /sn:0 {0}(1,1)(1,1){1}
wire w306;    //: /sn:0 {0}(1,1)(1,1){1}
wire w129;    //: /sn:0 {0}(1,1)(1,1){1}
wire w686;    //: /sn:0 {0}(1,1)(1,1){1}
wire w331;    //: /sn:0 {0}(1,1)(1,1){1}
wire w837;    //: /sn:0 {0}(1,1)(1,1){1}
wire w267;    //: /sn:0 {0}(1,1)(1,1){1}
wire w361;    //: /sn:0 {0}(1,1)(1,1){1}
wire w259;    //: /sn:0 {0}(1,1)(1,1){1}
wire w537;    //: /sn:0 {0}(1,1)(1,1){1}
wire w767;    //: /sn:0 {0}(1,1)(1,1){1}
wire w396;    //: /sn:0 {0}(1,1)(1,1){1}
wire w340;    //: /sn:0 {0}(1,1)(1,1){1}
wire w333;    //: /sn:0 {0}(1,1)(1,1){1}
wire w21;    //: /sn:0 {0}(1,1)(1,1){1}
wire w170;    //: /sn:0 {0}(1,1)(1,1){1}
wire w230;    //: /sn:0 {0}(1,1)(1,1){1}
wire w600;    //: /sn:0 {0}(1,1)(1,1){1}
wire w538;    //: /sn:0 {0}(1,1)(1,1){1}
wire w358;    //: /sn:0 {0}(1,1)(1,1){1}
wire w890;    //: /sn:0 {0}(1,1)(1,1){1}
wire w922;    //: /sn:0 {0}(1,1)(1,1){1}
wire w415;    //: /sn:0 {0}(1,1)(1,1){1}
wire w256;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1;    //: /sn:0 {0}(1,1)(1,1){1}
wire w674;    //: /sn:0 {0}(1,1)(1,1){1}
wire w776;    //: /sn:0 {0}(1,1)(1,1){1}
wire w409;    //: /sn:0 {0}(1,1)(1,1){1}
wire w241;    //: /sn:0 {0}(1,1)(1,1){1}
wire w941;    //: /sn:0 {0}(1,1)(1,1){1}
wire w584;    //: /sn:0 {0}(1,1)(1,1){1}
wire w655;    //: /sn:0 {0}(1,1)(1,1){1}
wire w98;    //: /sn:0 {0}(1,1)(1,1){1}
wire w116;    //: /sn:0 {0}(1,1)(1,1){1}
wire w798;    //: /sn:0 {0}(1,1)(1,1){1}
wire w338;    //: /sn:0 {0}(1,1)(1,1){1}
wire w869;    //: /sn:0 {0}(1,1)(1,1){1}
wire w198;    //: /sn:0 {0}(1,1)(1,1){1}
wire w702;    //: /sn:0 {0}(1,1)(1,1){1}
wire w11;    //: /sn:0 {0}(1,1)(1,1){1}
wire w137;    //: /sn:0 {0}(1,1)(1,1){1}
wire w193;    //: /sn:0 {0}(1,1)(1,1){1}
wire w611;    //: /sn:0 {0}(1,1)(1,1){1}
wire w717;    //: /sn:0 {0}(1,1)(1,1){1}
wire w848;    //: /sn:0 {0}(1,1)(1,1){1}
wire w923;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1003;    //: /sn:0 {0}(1,1)(1,1){1}
wire w13;    //: /sn:0 {0}(1,1)(1,1){1}
wire w208;    //: /sn:0 {0}(1,1)(1,1){1}
wire w410;    //: /sn:0 {0}(1,1)(1,1){1}
wire w131;    //: /sn:0 {0}(1,1)(1,1){1}
wire w471;    //: /sn:0 {0}(1,1)(1,1){1}
wire w823;    //: /sn:0 {0}(1,1)(1,1){1}
wire w390;    //: /sn:0 {0}(1,1)(1,1){1}
wire w278;    //: /sn:0 {0}(1,1)(1,1){1}
wire w737;    //: /sn:0 {0}(1,1)(1,1){1}
wire w341;    //: /sn:0 {0}(1,1)(1,1){1}
wire w160;    //: /sn:0 {0}(1,1)(1,1){1}
wire w704;    //: /sn:0 {0}(1,1)(1,1){1}
wire w392;    //: /sn:0 {0}(1,1)(1,1){1}
wire w526;    //: /sn:0 {0}(1,1)(1,1){1}
wire w566;    //: /sn:0 {0}(1,1)(1,1){1}
wire w151;    //: /sn:0 {0}(1,1)(1,1){1}
wire w657;    //: /sn:0 {0}(1,1)(1,1){1}
wire w692;    //: /sn:0 {0}(1,1)(1,1){1}
wire w397;    //: /sn:0 {0}(1,1)(1,1){1}
wire w582;    //: /sn:0 {0}(1,1)(1,1){1}
wire w368;    //: /sn:0 {0}(1,1)(1,1){1}
wire w104;    //: /sn:0 {0}(1,1)(1,1){1}
wire w111;    //: /sn:0 {0}(1,1)(1,1){1}
wire w171;    //: /sn:0 {0}(1,1)(1,1){1}
wire w622;    //: /sn:0 {0}(1,1)(1,1){1}
wire w641;    //: /sn:0 {0}(1,1)(1,1){1}
wire w237;    //: /sn:0 {0}(1,1)(1,1){1}
wire w67;    //: /sn:0 {0}(1,1)(1,1){1}
wire w936;    //: /sn:0 {0}(1,1)(1,1){1}
wire w448;    //: /sn:0 {0}(1,1)(1,1){1}
wire w607;    //: /sn:0 {0}(1,1)(1,1){1}
wire w621;    //: /sn:0 {0}(1,1)(1,1){1}
wire w797;    //: /sn:0 {0}(1,1)(1,1){1}
wire w920;    //: /sn:0 {0}(1,1)(1,1){1}
wire w369;    //: /sn:0 {0}(1,1)(1,1){1}
wire w298;    //: /sn:0 {0}(1,1)(1,1){1}
wire w108;    //: /sn:0 {0}(1,1)(1,1){1}
wire w985;    //: /sn:0 {0}(1,1)(1,1){1}
wire w223;    //: /sn:0 {0}(1,1)(1,1){1}
wire w827;    //: /sn:0 {0}(1,1)(1,1){1}
wire w951;    //: /sn:0 {0}(1,1)(1,1){1}
wire w8;    //: /sn:0 {0}(1,1)(1,1){1}
wire w573;    //: /sn:0 {0}(1,1)(1,1){1}
wire w814;    //: /sn:0 {0}(1,1)(1,1){1}
wire w202;    //: /sn:0 {0}(1,1)(1,1){1}
wire w669;    //: /sn:0 {0}(1,1)(1,1){1}
wire w84;    //: /sn:0 {0}(1,1)(1,1){1}
wire w755;    //: /sn:0 {0}(1,1)(1,1){1}
wire w821;    //: /sn:0 {0}(1,1)(1,1){1}
wire w850;    //: /sn:0 {0}(1,1)(1,1){1}
wire w362;    //: /sn:0 {0}(1,1)(1,1){1}
wire w351;    //: /sn:0 {0}(1,1)(1,1){1}
wire w315;    //: /sn:0 {0}(1,1)(1,1){1}
wire w274;    //: /sn:0 {0}(1,1)(1,1){1}
wire w458;    //: /sn:0 {0}(1,1)(1,1){1}
wire w695;    //: /sn:0 {0}(1,1)(1,1){1}
wire w347;    //: /sn:0 {0}(1,1)(1,1){1}
wire w52;    //: /sn:0 {0}(1,1)(1,1){1}
wire w461;    //: /sn:0 {0}(1,1)(1,1){1}
wire w510;    //: /sn:0 {0}(1,1)(1,1){1}
wire w596;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1011;    //: /sn:0 {0}(1,1)(1,1){1}
wire w696;    //: /sn:0 {0}(1,1)(1,1){1}
wire w913;    //: /sn:0 {0}(1,1)(1,1){1}
wire w416;    //: /sn:0 {0}(1,1)(1,1){1}
wire w406;    //: /sn:0 {0}(1,1)(1,1){1}
wire w329;    //: /sn:0 {0}(1,1)(1,1){1}
wire w550;    //: /sn:0 {0}(1,1)(1,1){1}
wire w683;    //: /sn:0 {0}(1,1)(1,1){1}
wire w69;    //: /sn:0 {0}(1,1)(1,1){1}
wire w290;    //: /sn:0 {0}(1,1)(1,1){1}
wire w271;    //: /sn:0 {0}(1,1)(1,1){1}
wire w66;    //: /sn:0 {0}(1,1)(1,1){1}
wire w177;    //: /sn:0 {0}(1,1)(1,1){1}
wire w891;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1020;    //: /sn:0 {0}(1,1)(1,1){1}
wire w234;    //: /sn:0 {0}(1,1)(1,1){1}
wire w761;    //: /sn:0 {0}(1,1)(1,1){1}
wire w835;    //: /sn:0 {0}(1,1)(1,1){1}
wire w326;    //: /sn:0 {0}(1,1)(1,1){1}
wire w323;    //: /sn:0 {0}(1,1)(1,1){1}
wire w87;    //: /sn:0 {0}(1,1)(1,1){1}
wire w534;    //: /sn:0 {0}(1,1)(1,1){1}
wire w829;    //: /sn:0 {0}(1,1)(1,1){1}
wire w375;    //: /sn:0 {0}(1,1)(1,1){1}
wire w321;    //: /sn:0 {0}(1,1)(1,1){1}
wire w307;    //: /sn:0 {0}(1,1)(1,1){1}
wire w28;    //: /sn:0 {0}(1,1)(1,1){1}
wire w130;    //: /sn:0 {0}(1,1)(1,1){1}
wire w698;    //: /sn:0 {0}(1,1)(1,1){1}
wire w385;    //: /sn:0 {0}(1,1)(1,1){1}
wire w833;    //: /sn:0 {0}(1,1)(1,1){1}
wire w343;    //: /sn:0 {0}(1,1)(1,1){1}
wire w377;    //: /sn:0 {0}(1,1)(1,1){1}
wire w25;    //: /sn:0 {0}(1,1)(1,1){1}
wire w925;    //: /sn:0 {0}(1,1)(1,1){1}
wire w681;    //: /sn:0 {0}(1,1)(1,1){1}
wire w121;    //: /sn:0 {0}(1,1)(1,1){1}
wire w488;    //: /sn:0 {0}(1,1)(1,1){1}
wire w470;    //: /sn:0 {0}(1,1)(1,1){1}
wire w736;    //: /sn:0 {0}(1,1)(1,1){1}
wire w995;    //: /sn:0 {0}(1,1)(1,1){1}
wire w355;    //: /sn:0 {0}(1,1)(1,1){1}
wire w912;    //: /sn:0 {0}(1,1)(1,1){1}
wire w248;    //: /sn:0 {0}(1,1)(1,1){1}
wire w581;    //: /sn:0 {0}(1,1)(1,1){1}
wire w831;    //: /sn:0 {0}(1,1)(1,1){1}
wire w49;    //: /sn:0 {0}(1,1)(1,1){1}
wire w139;    //: /sn:0 {0}(1,1)(1,1){1}
wire w418;    //: /sn:0 {0}(1,1)(1,1){1}
wire w680;    //: /sn:0 {0}(1,1)(1,1){1}
wire w861;    //: /sn:0 {0}(1,1)(1,1){1}
wire w268;    //: /sn:0 {0}(1,1)(1,1){1}
wire w580;    //: /sn:0 {0}(1,1)(1,1){1}
wire w682;    //: /sn:0 {0}(1,1)(1,1){1}
wire w973;    //: /sn:0 {0}(1,1)(1,1){1}
wire w191;    //: /sn:0 {0}(1,1)(1,1){1}
wire w597;    //: /sn:0 {0}(1,1)(1,1){1}
wire w684;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1012;    //: /sn:0 {0}(1,1)(1,1){1}
wire w107;    //: /sn:0 {0}(1,1)(1,1){1}
wire w805;    //: /sn:0 {0}(1,1)(1,1){1}
wire w436;    //: /sn:0 {0}(1,1)(1,1){1}
wire w536;    //: /sn:0 {0}(1,1)(1,1){1}
wire w279;    //: /sn:0 {0}(1,1)(1,1){1}
wire w232;    //: /sn:0 {0}(1,1)(1,1){1}
wire w430;    //: /sn:0 {0}(1,1)(1,1){1}
wire w563;    //: /sn:0 {0}(1,1)(1,1){1}
wire w134;    //: /sn:0 {0}(1,1)(1,1){1}
wire w733;    //: /sn:0 {0}(1,1)(1,1){1}
wire w880;    //: /sn:0 {0}(1,1)(1,1){1}
wire w179;    //: /sn:0 {0}(1,1)(1,1){1}
wire w528;    //: /sn:0 {0}(1,1)(1,1){1}
wire w452;    //: /sn:0 {0}(1,1)(1,1){1}
wire w846;    //: /sn:0 {0}(1,1)(1,1){1}
wire w841;    //: /sn:0 {0}(1,1)(1,1){1}
wire w424;    //: /sn:0 {0}(1,1)(1,1){1}
wire w204;    //: /sn:0 {0}(1,1)(1,1){1}
wire w483;    //: /sn:0 {0}(1,1)(1,1){1}
wire w894;    //: /sn:0 {0}(1,1)(1,1){1}
wire w990;    //: /sn:0 {0}(1,1)(1,1){1}
wire w501;    //: /sn:0 {0}(1,1)(1,1){1}
wire w504;    //: /sn:0 {0}(1,1)(1,1){1}
wire w729;    //: /sn:0 {0}(1,1)(1,1){1}
wire w759;    //: /sn:0 {0}(1,1)(1,1){1}
wire w311;    //: /sn:0 {0}(1,1)(1,1){1}
wire w156;    //: /sn:0 {0}(1,1)(1,1){1}
wire w524;    //: /sn:0 {0}(1,1)(1,1){1}
wire w335;    //: /sn:0 {0}(1,1)(1,1){1}
wire w532;    //: /sn:0 {0}(1,1)(1,1){1}
wire w242;    //: /sn:0 {0}(1,1)(1,1){1}
wire w491;    //: /sn:0 {0}(1,1)(1,1){1}
wire w280;    //: /sn:0 {0}(1,1)(1,1){1}
wire w903;    //: /sn:0 {0}(1,1)(1,1){1}
wire w933;    //: /sn:0 {0}(1,1)(1,1){1}
wire w974;    //: /sn:0 {0}(1,1)(1,1){1}
wire w35;    //: /sn:0 {0}(1,1)(1,1){1}
wire w91;    //: /sn:0 {0}(1,1)(1,1){1}
wire w477;    //: /sn:0 {0}(1,1)(1,1){1}
wire w591;    //: /sn:0 {0}(1,1)(1,1){1}
wire w163;    //: /sn:0 {0}(1,1)(1,1){1}
wire w765;    //: /sn:0 {0}(1,1)(1,1){1}
wire w332;    //: /sn:0 {0}(1,1)(1,1){1}
wire w144;    //: /sn:0 {0}(1,1)(1,1){1}
wire w557;    //: /sn:0 {0}(1,1)(1,1){1}
wire w716;    //: /sn:0 {0}(1,1)(1,1){1}
wire w554;    //: /sn:0 {0}(1,1)(1,1){1}
wire w659;    //: /sn:0 {0}(1,1)(1,1){1}
wire w228;    //: /sn:0 {0}(1,1)(1,1){1}
wire w12;    //: /sn:0 {0}(1,1)(1,1){1}
wire w543;    //: /sn:0 {0}(1,1)(1,1){1}
wire w309;    //: /sn:0 {0}(1,1)(1,1){1}
wire w365;    //: /sn:0 {0}(1,1)(1,1){1}
wire w583;    //: /sn:0 {0}(1,1)(1,1){1}
wire w257;    //: /sn:0 {0}(1,1)(1,1){1}
wire w27;    //: /sn:0 {0}(1,1)(1,1){1}
wire w455;    //: /sn:0 {0}(1,1)(1,1){1}
wire w549;    //: /sn:0 {0}(1,1)(1,1){1}
wire w914;    //: /sn:0 {0}(1,1)(1,1){1}
wire w468;    //: /sn:0 {0}(1,1)(1,1){1}
wire w870;    //: /sn:0 {0}(1,1)(1,1){1}
wire w489;    //: /sn:0 {0}(1,1)(1,1){1}
wire w921;    //: /sn:0 {0}(1,1)(1,1){1}
wire w378;    //: /sn:0 {0}(1,1)(1,1){1}
wire w281;    //: /sn:0 {0}(1,1)(1,1){1}
wire w412;    //: /sn:0 {0}(1,1)(1,1){1}
wire w966;    //: /sn:0 {0}(1,1)(1,1){1}
wire w637;    //: /sn:0 {0}(1,1)(1,1){1}
wire w516;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1023;    //: /sn:0 {0}(1,1)(1,1){1}
wire w414;    //: /sn:0 {0}(1,1)(1,1){1}
wire w539;    //: /sn:0 {0}(1,1)(1,1){1}
wire w838;    //: /sn:0 {0}(1,1)(1,1){1}
wire w63;    //: /sn:0 {0}(1,1)(1,1){1}
wire w159;    //: /sn:0 {0}(1,1)(1,1){1}
wire w627;    //: /sn:0 {0}(1,1)(1,1){1}
wire w236;    //: /sn:0 {0}(1,1)(1,1){1}
wire w76;    //: /sn:0 {0}(1,1)(1,1){1}
wire w545;    //: /sn:0 {0}(1,1)(1,1){1}
wire w594;    //: /sn:0 {0}(1,1)(1,1){1}
wire w434;    //: /sn:0 {0}(1,1)(1,1){1}
wire w199;    //: /sn:0 {0}(1,1)(1,1){1}
wire w712;    //: /sn:0 {0}(1,1)(1,1){1}
wire w249;    //: /sn:0 {0}(1,1)(1,1){1}
wire w968;    //: /sn:0 {0}(1,1)(1,1){1}
wire w551;    //: /sn:0 {0}(1,1)(1,1){1}
wire w884;    //: /sn:0 {0}(1,1)(1,1){1}
wire w658;    //: /sn:0 {0}(1,1)(1,1){1}
wire w840;    //: /sn:0 {0}(1,1)(1,1){1}
wire w328;    //: /sn:0 {0}(1,1)(1,1){1}
wire w260;    //: /sn:0 {0}(1,1)(1,1){1}
wire w889;    //: /sn:0 {0}(1,1)(1,1){1}
wire w403;    //: /sn:0 {0}(1,1)(1,1){1}
wire w310;    //: /sn:0 {0}(1,1)(1,1){1}
wire w541;    //: /sn:0 {0}(1,1)(1,1){1}
wire w253;    //: /sn:0 {0}(1,1)(1,1){1}
wire w522;    //: /sn:0 {0}(1,1)(1,1){1}
wire w786;    //: /sn:0 {0}(1,1)(1,1){1}
wire w371;    //: /sn:0 {0}(1,1)(1,1){1}
wire w590;    //: /sn:0 {0}(1,1)(1,1){1}
wire w656;    //: /sn:0 {0}(1,1)(1,1){1}
wire w739;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1018;    //: /sn:0 {0}(1,1)(1,1){1}
wire w123;    //: /sn:0 {0}(1,1)(1,1){1}
wire w993;    //: /sn:0 {0}(1,1)(1,1){1}
wire w969;    //: /sn:0 {0}(1,1)(1,1){1}
wire w427;    //: /sn:0 {0}(1,1)(1,1){1}
wire w295;    //: /sn:0 {0}(1,1)(1,1){1}
wire w185;    //: /sn:0 {0}(1,1)(1,1){1}
wire w568;    //: /sn:0 {0}(1,1)(1,1){1}
wire w807;    //: /sn:0 {0}(1,1)(1,1){1}
wire w924;    //: /sn:0 {0}(1,1)(1,1){1}
wire w319;    //: /sn:0 {0}(1,1)(1,1){1}
wire w930;    //: /sn:0 {0}(1,1)(1,1){1}
wire w293;    //: /sn:0 {0}(1,1)(1,1){1}
wire w70;    //: /sn:0 {0}(1,1)(1,1){1}
wire w766;    //: /sn:0 {0}(1,1)(1,1){1}
wire w906;    //: /sn:0 {0}(1,1)(1,1){1}
wire w497;    //: /sn:0 {0}(1,1)(1,1){1}
wire w88;    //: /sn:0 {0}(1,1)(1,1){1}
wire w565;    //: /sn:0 {0}(1,1)(1,1){1}
wire w47;    //: /sn:0 {0}(1,1)(1,1){1}
wire w642;    //: /sn:0 {0}(1,1)(1,1){1}
wire w862;    //: /sn:0 {0}(1,1)(1,1){1}
wire w806;    //: /sn:0 {0}(1,1)(1,1){1}
wire w512;    //: /sn:0 {0}(1,1)(1,1){1}
//: enddecls

  //: IN g4 (E4) @(1,1) /sn:0 /w:[ 0 ]
  //: IN g8 (E8) @(1,1) /sn:0 /w:[ 0 ]
  //: IN g13 (E13) @(1,1) /sn:0 /w:[ 0 ]
  //: OUT g37 (S5) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g55 (S23) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g58 (S26) @(1,1) /sn:0 /w:[ 1 ]
  assign S16 = {w1008, w976, w944, w912, w880, w848, w816, w784, w752, w720, w688, w656, w624, w592, w560, w528, w496, w464, w432, w400, w368, w336, w304, w272, w240, w208, w176, w144, w112, w80, w48, w16}; //: CONCAT g112  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign {w415, w414, w413, w412, w411, w410, w409, w408, w407, w406, w405, w404, w403, w402, w401, w400, w399, w398, w397, w396, w395, w394, w393, w392, w391, w390, w389, w388, w387, w386, w385, w384} = E12; //: CONCAT g76  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S15 = {w1007, w975, w943, w911, w879, w847, w815, w783, w751, w719, w687, w655, w623, w591, w559, w527, w495, w463, w431, w399, w367, w335, w303, w271, w239, w207, w175, w143, w111, w79, w47, w15}; //: CONCAT g111  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g1 (E1) @(1,1) /sn:0 /w:[ 0 ]
  assign {w31, w30, w29, w28, w27, w26, w25, w24, w23, w22, w21, w20, w19, w18, w17, w16, w15, w14, w13, w12, w11, w10, w9, w8, w7, w6, w5, w4, w3, w2, w1, w0} = E0; //: CONCAT g64  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: IN g11 (E11) @(1,1) /sn:0 /w:[ 0 ]
  assign S25 = {w1017, w985, w953, w921, w889, w857, w825, w793, w761, w729, w697, w665, w633, w601, w569, w537, w505, w473, w441, w409, w377, w345, w313, w281, w249, w217, w185, w153, w121, w89, w57, w25}; //: CONCAT g121  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g28 (E28) @(1,1) /sn:0 /w:[ 0 ]
  //: OUT g50 (S18) @(1,1) /sn:0 /w:[ 1 ]
  assign S17 = {w1009, w977, w945, w913, w881, w849, w817, w785, w753, w721, w689, w657, w625, w593, w561, w529, w497, w465, w433, w401, w369, w337, w305, w273, w241, w209, w177, w145, w113, w81, w49, w17}; //: CONCAT g113  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g19 (E19) @(1,1) /sn:0 /w:[ 0 ]
  assign S19 = {w1011, w979, w947, w915, w883, w851, w819, w787, w755, w723, w691, w659, w627, w595, w563, w531, w499, w467, w435, w403, w371, w339, w307, w275, w243, w211, w179, w147, w115, w83, w51, w19}; //: CONCAT g115  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g6 (E6) @(1,1) /sn:0 /w:[ 0 ]
  //: OUT g38 (S6) @(1,1) /sn:0 /w:[ 1 ]
  assign {w383, w382, w381, w380, w379, w378, w377, w376, w375, w374, w373, w372, w371, w370, w369, w368, w367, w366, w365, w364, w363, w362, w361, w360, w359, w358, w357, w356, w355, w354, w353, w352} = E11; //: CONCAT g75  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: IN g7 (E7) @(1,1) /sn:0 /w:[ 0 ]
  //: OUT g53 (S21) @(1,1) /sn:0 /w:[ 1 ]
  //: IN g20 (E20) @(1,1) /sn:0 /w:[ 0 ]
  //: IN g31 (E31) @(1,1) /sn:0 /w:[ 0 ]
  assign S28 = {w1020, w988, w956, w924, w892, w860, w828, w796, w764, w732, w700, w668, w636, w604, w572, w540, w508, w476, w444, w412, w380, w348, w316, w284, w252, w220, w188, w156, w124, w92, w60, w28}; //: CONCAT g124  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign {w159, w158, w157, w156, w155, w154, w153, w152, w151, w150, w149, w148, w147, w146, w145, w144, w143, w142, w141, w140, w139, w138, w137, w136, w135, w134, w133, w132, w131, w130, w129, w128} = E4; //: CONCAT g68  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: OUT g39 (S7) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g48 (S16) @(1,1) /sn:0 /w:[ 1 ]
  //: IN g17 (E17) @(1,1) /sn:0 /w:[ 0 ]
  //: IN g25 (E25) @(1,1) /sn:0 /w:[ 0 ]
  //: IN g29 (E29) @(1,1) /sn:0 /w:[ 0 ]
  assign S10 = {w1002, w970, w938, w906, w874, w842, w810, w778, w746, w714, w682, w650, w618, w586, w554, w522, w490, w458, w426, w394, w362, w330, w298, w266, w234, w202, w170, w138, w106, w74, w42, w10}; //: CONCAT g106  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S11 = {w1003, w971, w939, w907, w875, w843, w811, w779, w747, w715, w683, w651, w619, w587, w555, w523, w491, w459, w427, w395, w363, w331, w299, w267, w235, w203, w171, w139, w107, w75, w43, w11}; //: CONCAT g107  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g52 (S20) @(1,1) /sn:0 /w:[ 1 ]
  assign {w639, w638, w637, w636, w635, w634, w633, w632, w631, w630, w629, w628, w627, w626, w625, w624, w623, w622, w621, w620, w619, w618, w617, w616, w615, w614, w613, w612, w611, w610, w609, w608} = E19; //: CONCAT g83  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S4 = {w996, w964, w932, w900, w868, w836, w804, w772, w740, w708, w676, w644, w612, w580, w548, w516, w484, w452, w420, w388, w356, w324, w292, w260, w228, w196, w164, w132, w100, w68, w36, w4}; //: CONCAT g100  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g14 (E14) @(1,1) /sn:0 /w:[ 0 ]
  assign {w543, w542, w541, w540, w539, w538, w537, w536, w535, w534, w533, w532, w531, w530, w529, w528, w527, w526, w525, w524, w523, w522, w521, w520, w519, w518, w517, w516, w515, w514, w513, w512} = E16; //: CONCAT g80  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w991, w990, w989, w988, w987, w986, w985, w984, w983, w982, w981, w980, w979, w978, w977, w976, w975, w974, w973, w972, w971, w970, w969, w968, w967, w966, w965, w964, w963, w962, w961, w960} = E30; //: CONCAT g94  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: OUT g44 (S12) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g47 (S15) @(1,1) /sn:0 /w:[ 1 ]
  assign {w671, w670, w669, w668, w667, w666, w665, w664, w663, w662, w661, w660, w659, w658, w657, w656, w655, w654, w653, w652, w651, w650, w649, w648, w647, w646, w645, w644, w643, w642, w641, w640} = E20; //: CONCAT g84  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S9 = {w1001, w969, w937, w905, w873, w841, w809, w777, w745, w713, w681, w649, w617, w585, w553, w521, w489, w457, w425, w393, w361, w329, w297, w265, w233, w201, w169, w137, w105, w73, w41, w9}; //: CONCAT g105  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g21 (E21) @(1,1) /sn:0 /w:[ 0 ]
  //: IN g23 (E23) @(1,1) /sn:0 /w:[ 0 ]
  //: OUT g41 (S9) @(1,1) /sn:0 /w:[ 1 ]
  assign {w959, w958, w957, w956, w955, w954, w953, w952, w951, w950, w949, w948, w947, w946, w945, w944, w943, w942, w941, w940, w939, w938, w937, w936, w935, w934, w933, w932, w931, w930, w929, w928} = E29; //: CONCAT g93  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S20 = {w1012, w980, w948, w916, w884, w852, w820, w788, w756, w724, w692, w660, w628, w596, w564, w532, w500, w468, w436, w404, w372, w340, w308, w276, w244, w212, w180, w148, w116, w84, w52, w20}; //: CONCAT g116  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S27 = {w1019, w987, w955, w923, w891, w859, w827, w795, w763, w731, w699, w667, w635, w603, w571, w539, w507, w475, w443, w411, w379, w347, w315, w283, w251, w219, w187, w155, w123, w91, w59, w27}; //: CONCAT g123  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g40 (S8) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g54 (S22) @(1,1) /sn:0 /w:[ 1 ]
  assign {w863, w862, w861, w860, w859, w858, w857, w856, w855, w854, w853, w852, w851, w850, w849, w848, w847, w846, w845, w844, w843, w842, w841, w840, w839, w838, w837, w836, w835, w834, w833, w832} = E26; //: CONCAT g90  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: IN g0 (E0) @(1,1) /sn:0 /w:[ 0 ]
  //: IN g26 (E26) @(1,1) /sn:0 /w:[ 0 ]
  //: OUT g46 (S14) @(1,1) /sn:0 /w:[ 1 ]
  assign {w607, w606, w605, w604, w603, w602, w601, w600, w599, w598, w597, w596, w595, w594, w593, w592, w591, w590, w589, w588, w587, w586, w585, w584, w583, w582, w581, w580, w579, w578, w577, w576} = E18; //: CONCAT g82  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: comment g128 @(185,85) /sn:0
  //: /line:"Este modulo esta generado automaticamente con un programa. Estan todos los cables en el mismo punto por eso no se ven."
  //: /line:"Este modulo es para hcaer las conbinaciones de cables de um multiplexor."
  //: /end
  assign {w895, w894, w893, w892, w891, w890, w889, w888, w887, w886, w885, w884, w883, w882, w881, w880, w879, w878, w877, w876, w875, w874, w873, w872, w871, w870, w869, w868, w867, w866, w865, w864} = E27; //: CONCAT g91  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: OUT g33 (S1) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g49 (S17) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g61 (S29) @(1,1) /sn:0 /w:[ 1 ]
  assign {w735, w734, w733, w732, w731, w730, w729, w728, w727, w726, w725, w724, w723, w722, w721, w720, w719, w718, w717, w716, w715, w714, w713, w712, w711, w710, w709, w708, w707, w706, w705, w704} = E22; //: CONCAT g86  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: IN g3 (E3) @(1,1) /sn:0 /w:[ 0 ]
  //: OUT g34 (S2) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g51 (S19) @(1,1) /sn:0 /w:[ 1 ]
  assign {w831, w830, w829, w828, w827, w826, w825, w824, w823, w822, w821, w820, w819, w818, w817, w816, w815, w814, w813, w812, w811, w810, w809, w808, w807, w806, w805, w804, w803, w802, w801, w800} = E25; //: CONCAT g89  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w63, w62, w61, w60, w59, w58, w57, w56, w55, w54, w53, w52, w51, w50, w49, w48, w47, w46, w45, w44, w43, w42, w41, w40, w39, w38, w37, w36, w35, w34, w33, w32} = E1; //: CONCAT g65  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w447, w446, w445, w444, w443, w442, w441, w440, w439, w438, w437, w436, w435, w434, w433, w432, w431, w430, w429, w428, w427, w426, w425, w424, w423, w422, w421, w420, w419, w418, w417, w416} = E13; //: CONCAT g77  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S14 = {w1006, w974, w942, w910, w878, w846, w814, w782, w750, w718, w686, w654, w622, w590, w558, w526, w494, w462, w430, w398, w366, w334, w302, w270, w238, w206, w174, w142, w110, w78, w46, w14}; //: CONCAT g110  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g2 (E2) @(1,1) /sn:0 /w:[ 0 ]
  //: OUT g59 (S27) @(1,1) /sn:0 /w:[ 1 ]
  assign {w287, w286, w285, w284, w283, w282, w281, w280, w279, w278, w277, w276, w275, w274, w273, w272, w271, w270, w269, w268, w267, w266, w265, w264, w263, w262, w261, w260, w259, w258, w257, w256} = E8; //: CONCAT g72  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S2 = {w994, w962, w930, w898, w866, w834, w802, w770, w738, w706, w674, w642, w610, w578, w546, w514, w482, w450, w418, w386, w354, w322, w290, w258, w226, w194, w162, w130, w98, w66, w34, w2}; //: CONCAT g98  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S3 = {w995, w963, w931, w899, w867, w835, w803, w771, w739, w707, w675, w643, w611, w579, w547, w515, w483, w451, w419, w387, w355, w323, w291, w259, w227, w195, w163, w131, w99, w67, w35, w3}; //: CONCAT g99  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S0 = {w992, w960, w928, w896, w864, w832, w800, w768, w736, w704, w672, w640, w608, w576, w544, w512, w480, w448, w416, w384, w352, w320, w288, w256, w224, w192, w160, w128, w96, w64, w32, w0}; //: CONCAT g96  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g16 (E16) @(1,1) /sn:0 /w:[ 0 ]
  assign S7 = {w999, w967, w935, w903, w871, w839, w807, w775, w743, w711, w679, w647, w615, w583, w551, w519, w487, w455, w423, w391, w359, w327, w295, w263, w231, w199, w167, w135, w103, w71, w39, w7}; //: CONCAT g103  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S26 = {w1018, w986, w954, w922, w890, w858, w826, w794, w762, w730, w698, w666, w634, w602, w570, w538, w506, w474, w442, w410, w378, w346, w314, w282, w250, w218, w186, w154, w122, w90, w58, w26}; //: CONCAT g122  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign {w479, w478, w477, w476, w475, w474, w473, w472, w471, w470, w469, w468, w467, w466, w465, w464, w463, w462, w461, w460, w459, w458, w457, w456, w455, w454, w453, w452, w451, w450, w449, w448} = E14; //: CONCAT g78  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w767, w766, w765, w764, w763, w762, w761, w760, w759, w758, w757, w756, w755, w754, w753, w752, w751, w750, w749, w748, w747, w746, w745, w744, w743, w742, w741, w740, w739, w738, w737, w736} = E23; //: CONCAT g87  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: IN g10 (E10) @(1,1) /sn:0 /w:[ 0 ]
  //: IN g27 (E27) @(1,1) /sn:0 /w:[ 0 ]
  //: OUT g32 (S0) @(1,1) /sn:0 /w:[ 1 ]
  assign S6 = {w998, w966, w934, w902, w870, w838, w806, w774, w742, w710, w678, w646, w614, w582, w550, w518, w486, w454, w422, w390, w358, w326, w294, w262, w230, w198, w166, w134, w102, w70, w38, w6}; //: CONCAT g102  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign {w191, w190, w189, w188, w187, w186, w185, w184, w183, w182, w181, w180, w179, w178, w177, w176, w175, w174, w173, w172, w171, w170, w169, w168, w167, w166, w165, w164, w163, w162, w161, w160} = E5; //: CONCAT g69  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S23 = {w1015, w983, w951, w919, w887, w855, w823, w791, w759, w727, w695, w663, w631, w599, w567, w535, w503, w471, w439, w407, w375, w343, w311, w279, w247, w215, w183, w151, w119, w87, w55, w23}; //: CONCAT g119  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g9 (E9) @(1,1) /sn:0 /w:[ 0 ]
  //: OUT g57 (S25) @(1,1) /sn:0 /w:[ 1 ]
  assign {w255, w254, w253, w252, w251, w250, w249, w248, w247, w246, w245, w244, w243, w242, w241, w240, w239, w238, w237, w236, w235, w234, w233, w232, w231, w230, w229, w228, w227, w226, w225, w224} = E7; //: CONCAT g71  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: IN g15 (E15) @(1,1) /sn:0 /w:[ 0 ]
  assign {w127, w126, w125, w124, w123, w122, w121, w120, w119, w118, w117, w116, w115, w114, w113, w112, w111, w110, w109, w108, w107, w106, w105, w104, w103, w102, w101, w100, w99, w98, w97, w96} = E3; //: CONCAT g67  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S31 = {w1023, w991, w959, w927, w895, w863, w831, w799, w767, w735, w703, w671, w639, w607, w575, w543, w511, w479, w447, w415, w383, w351, w319, w287, w255, w223, w191, w159, w127, w95, w63, w31}; //: CONCAT g127  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g43 (S11) @(1,1) /sn:0 /w:[ 1 ]
  assign {w319, w318, w317, w316, w315, w314, w313, w312, w311, w310, w309, w308, w307, w306, w305, w304, w303, w302, w301, w300, w299, w298, w297, w296, w295, w294, w293, w292, w291, w290, w289, w288} = E9; //: CONCAT g73  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w799, w798, w797, w796, w795, w794, w793, w792, w791, w790, w789, w788, w787, w786, w785, w784, w783, w782, w781, w780, w779, w778, w777, w776, w775, w774, w773, w772, w771, w770, w769, w768} = E24; //: CONCAT g88  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S8 = {w1000, w968, w936, w904, w872, w840, w808, w776, w744, w712, w680, w648, w616, w584, w552, w520, w488, w456, w424, w392, w360, w328, w296, w264, w232, w200, w168, w136, w104, w72, w40, w8}; //: CONCAT g104  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g62 (S30) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g42 (S10) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g63 (S31) @(1,1) /sn:0 /w:[ 1 ]
  assign {w351, w350, w349, w348, w347, w346, w345, w344, w343, w342, w341, w340, w339, w338, w337, w336, w335, w334, w333, w332, w331, w330, w329, w328, w327, w326, w325, w324, w323, w322, w321, w320} = E10; //: CONCAT g74  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S13 = {w1005, w973, w941, w909, w877, w845, w813, w781, w749, w717, w685, w653, w621, w589, w557, w525, w493, w461, w429, w397, w365, w333, w301, w269, w237, w205, w173, w141, w109, w77, w45, w13}; //: CONCAT g109  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g5 (E5) @(1,1) /sn:0 /w:[ 0 ]
  //: OUT g56 (S24) @(1,1) /sn:0 /w:[ 1 ]
  assign {w511, w510, w509, w508, w507, w506, w505, w504, w503, w502, w501, w500, w499, w498, w497, w496, w495, w494, w493, w492, w491, w490, w489, w488, w487, w486, w485, w484, w483, w482, w481, w480} = E15; //: CONCAT g79  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w1023, w1022, w1021, w1020, w1019, w1018, w1017, w1016, w1015, w1014, w1013, w1012, w1011, w1010, w1009, w1008, w1007, w1006, w1005, w1004, w1003, w1002, w1001, w1000, w999, w998, w997, w996, w995, w994, w993, w992} = E31; //: CONCAT g95  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S21 = {w1013, w981, w949, w917, w885, w853, w821, w789, w757, w725, w693, w661, w629, w597, w565, w533, w501, w469, w437, w405, w373, w341, w309, w277, w245, w213, w181, w149, w117, w85, w53, w21}; //: CONCAT g117  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign {w703, w702, w701, w700, w699, w698, w697, w696, w695, w694, w693, w692, w691, w690, w689, w688, w687, w686, w685, w684, w683, w682, w681, w680, w679, w678, w677, w676, w675, w674, w673, w672} = E21; //: CONCAT g85  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w927, w926, w925, w924, w923, w922, w921, w920, w919, w918, w917, w916, w915, w914, w913, w912, w911, w910, w909, w908, w907, w906, w905, w904, w903, w902, w901, w900, w899, w898, w897, w896} = E28; //: CONCAT g92  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: IN g24 (E24) @(1,1) /sn:0 /w:[ 0 ]
  //: OUT g36 (S4) @(1,1) /sn:0 /w:[ 1 ]
  assign S29 = {w1021, w989, w957, w925, w893, w861, w829, w797, w765, w733, w701, w669, w637, w605, w573, w541, w509, w477, w445, w413, w381, w349, w317, w285, w253, w221, w189, w157, w125, w93, w61, w29}; //: CONCAT g125  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign {w575, w574, w573, w572, w571, w570, w569, w568, w567, w566, w565, w564, w563, w562, w561, w560, w559, w558, w557, w556, w555, w554, w553, w552, w551, w550, w549, w548, w547, w546, w545, w544} = E17; //: CONCAT g81  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S5 = {w997, w965, w933, w901, w869, w837, w805, w773, w741, w709, w677, w645, w613, w581, w549, w517, w485, w453, w421, w389, w357, w325, w293, w261, w229, w197, w165, w133, w101, w69, w37, w5}; //: CONCAT g101  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g60 (S28) @(1,1) /sn:0 /w:[ 1 ]
  assign {w223, w222, w221, w220, w219, w218, w217, w216, w215, w214, w213, w212, w211, w210, w209, w208, w207, w206, w205, w204, w203, w202, w201, w200, w199, w198, w197, w196, w195, w194, w193, w192} = E6; //: CONCAT g70  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S30 = {w1022, w990, w958, w926, w894, w862, w830, w798, w766, w734, w702, w670, w638, w606, w574, w542, w510, w478, w446, w414, w382, w350, w318, w286, w254, w222, w190, w158, w126, w94, w62, w30}; //: CONCAT g126  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g22 (E22) @(1,1) /sn:0 /w:[ 0 ]
  //: OUT g35 (S3) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g45 (S13) @(1,1) /sn:0 /w:[ 1 ]
  assign {w95, w94, w93, w92, w91, w90, w89, w88, w87, w86, w85, w84, w83, w82, w81, w80, w79, w78, w77, w76, w75, w74, w73, w72, w71, w70, w69, w68, w67, w66, w65, w64} = E2; //: CONCAT g66  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S1 = {w993, w961, w929, w897, w865, w833, w801, w769, w737, w705, w673, w641, w609, w577, w545, w513, w481, w449, w417, w385, w353, w321, w289, w257, w225, w193, w161, w129, w97, w65, w33, w1}; //: CONCAT g97  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S18 = {w1010, w978, w946, w914, w882, w850, w818, w786, w754, w722, w690, w658, w626, w594, w562, w530, w498, w466, w434, w402, w370, w338, w306, w274, w242, w210, w178, w146, w114, w82, w50, w18}; //: CONCAT g114  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S24 = {w1016, w984, w952, w920, w888, w856, w824, w792, w760, w728, w696, w664, w632, w600, w568, w536, w504, w472, w440, w408, w376, w344, w312, w280, w248, w216, w184, w152, w120, w88, w56, w24}; //: CONCAT g120  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g12 (E12) @(1,1) /sn:0 /w:[ 0 ]
  //: IN g18 (E18) @(1,1) /sn:0 /w:[ 0 ]
  assign S12 = {w1004, w972, w940, w908, w876, w844, w812, w780, w748, w716, w684, w652, w620, w588, w556, w524, w492, w460, w428, w396, w364, w332, w300, w268, w236, w204, w172, w140, w108, w76, w44, w12}; //: CONCAT g108  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g30 (E30) @(1,1) /sn:0 /w:[ 0 ]
  assign S22 = {w1014, w982, w950, w918, w886, w854, w822, w790, w758, w726, w694, w662, w630, w598, w566, w534, w502, w470, w438, w406, w374, w342, w310, w278, w246, w214, w182, w150, w118, w86, w54, w22}; //: CONCAT g118  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1

endmodule
//: /netlistEnd

//: /netlistBegin Memoria
module Memoria(Esc, W, Direc, Reloj, Leer);
//: interface  /sz:(81, 80) /bd:[ Ti0>W(38/81) Li0>Direc[31:0](19/80) Li1>Esc[31:0](50/80) Bi0>Reloj(39/81) Ro0<Leer[31:0](37/80) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [31:0] Direc;    //: /sn:0 {0}(#:97,329)(174,329)(174,330)(#:248,330){1}
output [31:0] Leer;    //: /sn:0 {0}(707,235)(#:633,235){1}
input [31:0] Esc;    //: /sn:0 {0}(#:425,283)(#:503,283){1}
input Reloj;    //: /sn:0 {0}(569,348)(569,315)(568,315)(568,311){1}
input W;    //: /sn:0 {0}(565,146)(565,197){1}
supply0 w9;    //: /sn:0 {0}(451,154)(451,145)(450,145)(450,135){1}
//: {2}(452,133)(461,133)(461,154){3}
//: {4}(450,131)(450,125)(441,125)(441,154){5}
//: {6}(448,133)(423,133){7}
//: {8}(421,135)(421,125)(431,125)(431,154){9}
//: {10}(419,133)(377,133)(377,149){11}
//: {12}(421,135)(421,154){13}
wire w6;    //: /sn:0 {0}(321,225)(254,225){1}
wire w32;    //: /sn:0 {0}(254,395)(269,395){1}
wire [31:0] w7;    //: /sn:0 {0}(#:633,270)(648,270){1}
wire w4;    //: /sn:0 {0}(269,175)(254,175){1}
wire w19;    //: /sn:0 {0}(254,265)(269,265){1}
wire w38;    //: /sn:0 {0}(254,455)(269,455){1}
wire [4:0] w0;    //: /sn:0 {0}(#:441,160)(441,236)(#:503,236){1}
wire w3;    //: /sn:0 {0}(254,205)(321,205){1}
wire w37;    //: /sn:0 {0}(254,445)(269,445){1}
wire w34;    //: /sn:0 {0}(254,415)(269,415){1}
wire w21;    //: /sn:0 {0}(254,285)(269,285){1}
wire w31;    //: /sn:0 {0}(254,385)(269,385){1}
wire w28;    //: /sn:0 {0}(254,355)(269,355){1}
wire w20;    //: /sn:0 {0}(254,275)(269,275){1}
wire w23;    //: /sn:0 {0}(254,305)(269,305){1}
wire w24;    //: /sn:0 {0}(254,315)(269,315){1}
wire w36;    //: /sn:0 {0}(254,435)(269,435){1}
wire w41;    //: /sn:0 {0}(254,485)(269,485){1}
wire w1;    //: /sn:0 {0}(269,185)(254,185){1}
wire w25;    //: /sn:0 {0}(254,325)(269,325){1}
wire w8;    //: /sn:0 {0}(254,235)(321,235){1}
wire w18;    //: /sn:0 {0}(254,255)(269,255){1}
wire w35;    //: /sn:0 {0}(254,425)(269,425){1}
wire w40;    //: /sn:0 {0}(254,475)(269,475){1}
wire w30;    //: /sn:0 {0}(254,375)(269,375){1}
wire w17;    //: /sn:0 {0}(254,245)(269,245){1}
wire w22;    //: /sn:0 {0}(254,295)(269,295){1}
wire [4:0] w2;    //: /sn:0 {0}(#:327,215)(383,215){1}
//: {2}(387,215)(#:503,215){3}
//: {4}(385,217)(385,261)(#:503,261){5}
wire w12;    //: /sn:0 {0}(254,195)(321,195){1}
wire w27;    //: /sn:0 {0}(254,345)(269,345){1}
wire w5;    //: /sn:0 {0}(321,215)(254,215){1}
wire w33;    //: /sn:0 {0}(254,405)(269,405){1}
wire w29;    //: /sn:0 {0}(254,365)(269,365){1}
wire w26;    //: /sn:0 {0}(254,335)(269,335){1}
wire w39;    //: /sn:0 {0}(254,465)(269,465){1}
//: enddecls

  //: IN g4 (Esc) @(423,283) /sn:0 /w:[ 0 ]
  //: GROUND g8 (w9) @(377,155) /sn:0 /w:[ 11 ]
  //: IN g3 (W) @(565,144) /sn:0 /R:3 /w:[ 0 ]
  //: IN g13 (Direc) @(95,329) /sn:0 /w:[ 0 ]
  //: IN g2 (Reloj) @(569,350) /sn:0 /R:1 /w:[ 0 ]
  //: comment g1 @(281,96) /sn:0
  //: /line:"Esto no esta echo como en los apuntes"
  //: /end
  assign w2 = {w8, w6, w5, w3, w12}; //: CONCAT g11  @(326,215) /sn:0 /w:[ 0 1 0 0 1 1 ] /dr:1 /tp:0 /drp:1
  //: joint g10 (w9) @(450, 133) /w:[ 2 4 6 1 ]
  //: joint g6 (w2) @(385, 215) /w:[ 2 -1 1 4 ]
  assign w0 = {w9, w9, w9, w9, w9}; //: CONCAT g7  @(441,159) /sn:0 /R:3 /w:[ 0 3 0 5 9 13 ] /dr:0 /tp:0 /drp:1
  //: joint g9 (w9) @(421, 133) /w:[ 7 8 10 12 ]
  //: OUT g5 (Leer) @(704,235) /sn:0 /w:[ 0 ]
  Banco32Reg g0 (.W(W), .RegLeer2(w0), .RegLeer1(w2), .RegEsc(w2), .Esc(Esc), .Reloj(Reloj), .Leer2(w7), .Leer1(Leer));   //: @(504, 198) /sz:(128, 112) /sn:0 /p:[ Ti0>1 Li0>1 Li1>3 Li2>5 Li3>1 Bi0>1 Ro0<0 Ro1<1 ]
  assign {w41, w40, w39, w38, w37, w36, w35, w34, w33, w32, w31, w30, w29, w28, w27, w26, w25, w24, w23, w22, w21, w20, w19, w18, w17, w8, w6, w5, w3, w12, w1, w4} = Direc; //: CONCAT g12  @(249,330) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 ] /dr:0 /tp:0 /drp:0

endmodule
//: /netlistEnd

//: /netlistBegin Desplazador2
module Desplazador2(Sa, E);
//: interface  /sz:(88, 40) /bd:[ Li0>E[31:0](16/40) Ro0<Sa[31:0](16/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output [31:0] Sa;    //: /sn:0 {0}(#:497,250)(497,335)(544,335){1}
supply0 w2;    //: /sn:0 {0}(642,244)(642,224)(650,224){1}
//: {2}(654,224)(721,224)(721,262){3}
//: {4}(652,226)(652,244){5}
input [31:0] E;    //: /sn:0 {0}(#:477,191)(477,77)(#:437,77){1}
wire w6;    //: /sn:0 {0}(582,244)(582,197){1}
wire w32;    //: /sn:0 {0}(322,197)(322,212){1}
wire w7;    //: /sn:0 {0}(572,244)(572,197){1}
wire w14;    //: /sn:0 {0}(502,244)(502,197){1}
wire w16;    //: /sn:0 {0}(482,244)(482,197){1}
wire w4;    //: /sn:0 {0}(602,197)(602,244){1}
wire w15;    //: /sn:0 {0}(492,244)(492,197){1}
wire w19;    //: /sn:0 {0}(452,244)(452,197){1}
wire w0;    //: /sn:0 {0}(632,244)(632,197){1}
wire w3;    //: /sn:0 {0}(612,244)(612,197){1}
wire w21;    //: /sn:0 {0}(432,244)(432,197){1}
wire w31;    //: /sn:0 {0}(332,197)(332,212){1}
wire w28;    //: /sn:0 {0}(362,244)(362,197){1}
wire w20;    //: /sn:0 {0}(442,244)(442,197){1}
wire w23;    //: /sn:0 {0}(412,244)(412,197){1}
wire w24;    //: /sn:0 {0}(402,244)(402,197){1}
wire w1;    //: /sn:0 {0}(622,244)(622,197){1}
wire w25;    //: /sn:0 {0}(392,197)(392,244){1}
wire w8;    //: /sn:0 {0}(562,244)(562,197){1}
wire w18;    //: /sn:0 {0}(462,244)(462,197){1}
wire w30;    //: /sn:0 {0}(342,244)(342,197){1}
wire w17;    //: /sn:0 {0}(472,244)(472,197){1}
wire w22;    //: /sn:0 {0}(422,244)(422,197){1}
wire w11;    //: /sn:0 {0}(532,244)(532,197){1}
wire w12;    //: /sn:0 {0}(522,244)(522,197){1}
wire w10;    //: /sn:0 {0}(542,244)(542,197){1}
wire w13;    //: /sn:0 {0}(512,244)(512,197){1}
wire w27;    //: /sn:0 {0}(372,244)(372,197){1}
wire w5;    //: /sn:0 {0}(592,244)(592,197){1}
wire w29;    //: /sn:0 {0}(352,197)(352,244){1}
wire w9;    //: /sn:0 {0}(552,244)(552,197){1}
wire w26;    //: /sn:0 {0}(382,244)(382,197){1}
//: enddecls

  //: GROUND g4 (w2) @(721,268) /sn:0 /w:[ 3 ]
  //: OUT g3 (Sa) @(541,335) /sn:0 /w:[ 1 ]
  assign Sa = {w30, w29, w28, w27, w26, w25, w24, w23, w22, w21, w20, w19, w18, w17, w16, w15, w14, w13, w12, w11, w10, w9, w8, w7, w6, w5, w4, w3, w1, w0, w2, w2}; //: CONCAT g2  @(497,249) /sn:0 /R:3 /w:[ 0 0 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 5 ] /dr:1 /tp:0 /drp:1
  //: IN g1 (E) @(435,77) /sn:0 /w:[ 1 ]
  //: joint g5 (w2) @(652, 224) /w:[ 2 -1 1 4 ]
  assign {w32, w31, w30, w29, w28, w27, w26, w25, w24, w23, w22, w21, w20, w19, w18, w17, w16, w15, w14, w13, w12, w11, w10, w9, w8, w7, w6, w5, w4, w3, w1, w0} = E; //: CONCAT g0  @(477,192) /sn:0 /R:1 /w:[ 0 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 1 1 0 ] /dr:0 /tp:0 /drp:0

endmodule
//: /netlistEnd

//: /netlistBegin FlipFlopD
module FlipFlopD(Reloj, nQ, Q, W, D);
//: interface  /sz:(40, 40) /bd:[ Li0>D(6/40) Li1>Reloj(29/40) Bi0>W(33/40) Ro0<Q(5/40) Ro1<nQ(19/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output nQ;    //: /sn:0 {0}(458,135)(536,135)(536,191)(551,191){1}
output Q;    //: /sn:0 {0}(458,116)(551,116)(551,109)(566,109){1}
input D;    //: /sn:0 {0}(47,98)(158,98)(158,110)(188,110){1}
input Reloj;    //: /sn:0 {0}(46,293)(81,293)(81,281)(96,281){1}
input W;    //: /sn:0 {0}(374,327)(374,265){1}
//: {2}(374,261)(374,237)(359,237)(359,224){3}
//: {4}(372,263)(169,263)(169,224){5}
wire w3;    //: /sn:0 {0}(280,127)(265,127){1}
wire w0;    //: /sn:0 {0}(112,281)(139,281)(139,293)(162,293){1}
//: {2}(166,293)(196,293)(196,281)(207,281){3}
//: {4}(164,291)(164,224){5}
wire w1;    //: /sn:0 {0}(167,203)(167,125)(188,125){1}
wire w2;    //: /sn:0 {0}(265,108)(362,108)(362,118)(381,118){1}
wire w5;    //: /sn:0 {0}(357,203)(357,133)(381,133){1}
wire w9;    //: /sn:0 {0}(354,224)(354,281)(223,281){1}
//: enddecls

  //: IN g8 (Reloj) @(44,293) /sn:0 /w:[ 0 ]
  _GGAND2 #(6) g4 (.I0(w0), .I1(W), .Z(w1));   //: @(167,213) /sn:0 /R:1 /w:[ 5 5 0 ]
  //: OUT g3 (nQ) @(548,191) /sn:0 /w:[ 1 ]
  //: joint g13 (w0) @(164, 293) /w:[ 2 4 1 -1 ]
  //: OUT g2 (Q) @(563,109) /sn:0 /w:[ 1 ]
  LatchD g1 (.C(w5), .D(w2), .nQ(nQ), .Q(Q));   //: @(382, 104) /sz:(75, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  //: joint g11 (W) @(374, 263) /w:[ -1 2 4 1 ]
  _GGNBUF #(2) g10 (.I(Reloj), .Z(w0));   //: @(102,281) /sn:0 /w:[ 1 0 ]
  _GGNBUF #(2) g6 (.I(w0), .Z(w9));   //: @(213,281) /sn:0 /w:[ 3 1 ]
  //: IN g9 (W) @(374,329) /sn:0 /R:1 /w:[ 0 ]
  //: IN g7 (D) @(45,98) /sn:0 /w:[ 0 ]
  _GGAND2 #(6) g5 (.I0(w9), .I1(W), .Z(w5));   //: @(357,213) /sn:0 /R:1 /w:[ 0 3 0 ]
  LatchD g0 (.C(w1), .D(D), .nQ(w3), .Q(w2));   //: @(189, 96) /sz:(75, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  //: comment g12 @(343,29) /sn:0
  //: /line:"Flanco ascendente"
  //: /end

endmodule
//: /netlistEnd

//: /netlistBegin LatchSR
module LatchSR(Q, C, S, R, nQ);
//: interface  /sz:(81, 64) /bd:[ Li0>C(28/64) Li1>R(46/64) Li2>S(11/64) Ro0<nQ(40/64) Ro1<Q(20/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output Q;    //: /sn:0 {0}(443,120)(505,120)(505,112)(521,112){1}
//: {2}(525,112)(563,112){3}
//: {4}(523,114)(523,227)(404,227)(404,242)(414,242){5}
output nQ;    //: /sn:0 {0}(435,245)(500,245){1}
//: {2}(504,245)(561,245){3}
//: {4}(502,243)(502,137)(412,137)(412,122)(422,122){5}
input R;    //: /sn:0 {0}(156,97)(304,97)(304,114)(319,114){1}
input C;    //: /sn:0 {0}(173,192)(258,192){1}
//: {2}(260,190)(260,119)(319,119){3}
//: {4}(260,194)(260,258)(307,258){5}
input S;    //: /sn:0 {0}(196,295)(292,295)(292,263)(307,263){1}
wire w2;    //: /sn:0 {0}(340,117)(422,117){1}
wire w5;    //: /sn:0 {0}(328,261)(399,261)(399,247)(414,247){1}
//: enddecls

  //: OUT g4 (Q) @(560,112) /sn:0 /w:[ 3 ]
  //: IN g8 (C) @(171,192) /sn:0 /w:[ 0 ]
  _GGNOR2 #(4) g3 (.I0(Q), .I1(w5), .Z(nQ));   //: @(425,245) /sn:0 /w:[ 5 1 0 ]
  _GGNOR2 #(4) g2 (.I0(w2), .I1(nQ), .Z(Q));   //: @(433,120) /sn:0 /w:[ 1 5 0 ]
  _GGAND2 #(6) g1 (.I0(C), .I1(S), .Z(w5));   //: @(318,261) /sn:0 /w:[ 5 1 0 ]
  //: joint g11 (Q) @(523, 112) /w:[ 2 -1 1 4 ]
  //: joint g10 (nQ) @(502, 245) /w:[ 2 4 1 -1 ]
  //: IN g6 (S) @(194,295) /sn:0 /w:[ 0 ]
  //: IN g7 (R) @(154,97) /sn:0 /w:[ 0 ]
  //: joint g9 (C) @(260, 192) /w:[ -1 2 1 4 ]
  //: OUT g5 (nQ) @(558,245) /sn:0 /w:[ 3 ]
  _GGAND2 #(6) g0 (.I0(R), .I1(C), .Z(w2));   //: @(330,117) /sn:0 /w:[ 1 3 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin Mux5
module Mux5(E, C, Sa);
//: interface  /sz:(40, 40) /bd:[ Ti0>C[4:0](19/40) Li0>E[31:0](17/40) Ro0<Sa(19/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output Sa;    //: /sn:0 {0}(1267,628)(1363,628){1}
input [4:0] C;    //: /sn:0 {0}(#:97,-21)(97,-71)(94,-71)(#:94,-106){1}
input [31:0] E;    //: /sn:0 {0}(#:-584,633)(-471,633)(-471,645)(#:-427,645){1}
wire w6;    //: /sn:0 {0}(245,1184)(117,1184)(117,1153){1}
//: {2}(119,1151)(129,1151)(129,1152)(246,1152){3}
//: {4}(117,1149)(117,1126){5}
//: {6}(119,1124)(129,1124)(129,1121)(247,1121){7}
//: {8}(117,1122)(117,1093){9}
//: {10}(119,1091)(183,1091)(183,1089)(248,1089){11}
//: {12}(117,1089)(117,1053){13}
//: {14}(119,1051)(183,1051)(183,1049)(248,1049){15}
//: {16}(117,1049)(117,1022){17}
//: {18}(119,1020)(129,1020)(129,1017)(249,1017){19}
//: {20}(117,1018)(117,990){21}
//: {22}(119,988)(184,988)(184,985)(250,985){23}
//: {24}(117,986)(117,957){25}
//: {26}(119,955)(129,955)(129,954)(251,954){27}
//: {28}(117,953)(117,887){29}
//: {30}(119,885)(129,885)(129,884)(248,884){31}
//: {32}(117,883)(117,854){33}
//: {34}(119,852)(128,852)(128,852)(248,852){35}
//: {36}(117,850)(117,825){37}
//: {38}(119,823)(184,823)(184,821)(250,821){39}
//: {40}(117,821)(117,793){41}
//: {42}(119,791)(185,791)(185,788)(251,788){43}
//: {44}(117,789)(117,754){45}
//: {46}(119,752)(129,752)(129,749)(251,749){47}
//: {48}(117,750)(117,719){49}
//: {50}(119,717)(125,717)(125,718)(248,718){51}
//: {52}(117,715)(117,689){53}
//: {54}(119,687)(129,687)(129,686)(253,686){55}
//: {56}(117,685)(117,649){57}
//: {58}(119,647)(129,647)(129,654)(254,654){59}
//: {60}(117,645)(117,588){61}
//: {62}(119,586)(129,586)(129,589)(253,589){63}
//: {64}(117,584)(117,558){65}
//: {66}(119,556)(129,556)(129,557)(254,557){67}
//: {68}(117,554)(117,529){69}
//: {70}(119,527)(129,527)(129,526)(255,526){71}
//: {72}(117,525)(117,498){73}
//: {74}(119,496)(187,496)(187,494)(256,494){75}
//: {76}(117,494)(117,456){77}
//: {78}(119,454)(129,454)(129,454)(256,454){79}
//: {80}(117,452)(117,428){81}
//: {82}(119,426)(129,426)(129,422)(257,422){83}
//: {84}(117,424)(117,395){85}
//: {86}(119,393)(188,393)(188,391)(258,391){87}
//: {88}(117,391)(117,361){89}
//: {90}(119,359)(129,359)(129,359)(259,359){91}
//: {92}(117,357)(117,294){93}
//: {94}(119,292)(128,292)(128,289)(255,289){95}
//: {96}(117,290)(117,261){97}
//: {98}(119,259)(188,259)(188,257)(257,257){99}
//: {100}(117,257)(117,230){101}
//: {102}(119,228)(188,228)(188,226)(258,226){103}
//: {104}(117,226)(117,195){105}
//: {106}(119,193)(129,193)(129,194)(259,194){107}
//: {108}(117,191)(117,158){109}
//: {110}(119,156)(196,156)(196,153)(257,153){111}
//: {112}(117,154)(117,125){113}
//: {114}(119,123)(201,123)(201,122)(271,122){115}
//: {116}(117,121)(117,94){117}
//: {118}(119,92)(139,92)(139,89)(266,89){119}
//: {120}(117,90)(117,64){121}
//: {122}(119,62)(129,62)(129,59)(262,59){123}
//: {124}(117,60)(117,-15){125}
wire w32;    //: /sn:0 {0}(251,979)(-134,979)(-134,1045)(-149,1045){1}
wire w7;    //: /sn:0 {0}(271,147)(69,147)(69,159)(-155,159){1}
wire S1;    //: /sn:0 {0}(403,158)(380,158)(380,101)(287,101){1}
wire w73;    //: /sn:0 {0}(946,677)(1122,677)(1122,651)(1246,651){1}
wire w45;    //: /sn:0 {0}(1246,566)(1206,566)(1206,481)(946,481){1}
wire w61;    //: /sn:0 {0}(946,554)(1161,554)(1161,596)(1246,596){1}
wire w60;    //: /sn:0 {0}(946,544)(1172,544)(1172,591)(1246,591){1}
wire w46;    //: /sn:0 {0}(946,491)(1201,491)(1201,571)(1246,571){1}
wire S25;    //: /sn:0 {0}(271,997)(517,997)(517,1033)(576,1033){1}
wire w16;    //: /sn:0 {0}(257,447)(-158,447)(-158,452)(-173,452){1}
wire w14;    //: /sn:0 {0}(259,384)(-158,384)(-158,432)(-173,432){1}
wire w15;    //: /sn:0 {0}(258,416)(-146,416)(-146,442)(-173,442){1}
wire S6;    //: /sn:0 {0}(278,269)(370,269)(370,208)(403,208){1}
wire w81;    //: /sn:0 {0}(946,771)(1200,771)(1200,691)(1246,691){1}
wire w19;    //: /sn:0 {0}(255,551)(-121,551)(-121,482)(-173,482){1}
wire S7;    //: /sn:0 {0}(276,301)(387,301)(387,218)(403,218){1}
wire w4;    //: /sn:0 {0}(246,1167)(15,1167)(15,1168)(5,1168){1}
//: {2}(3,1166)(3,1137){3}
//: {4}(5,1135)(15,1135)(15,1136)(247,1136){5}
//: {6}(3,1133)(3,1108){7}
//: {8}(5,1106)(126,1106)(126,1104)(248,1104){9}
//: {10}(3,1104)(3,1066){11}
//: {12}(5,1064)(15,1064)(15,1064)(248,1064){13}
//: {14}(3,1062)(3,1030){15}
//: {16}(5,1028)(15,1028)(15,1032)(249,1032){17}
//: {18}(3,1026)(3,1004){19}
//: {20}(5,1002)(15,1002)(15,1000)(250,1000){21}
//: {22}(3,1000)(3,971){23}
//: {24}(5,969)(15,969)(15,969)(251,969){25}
//: {26}(3,967)(3,902){27}
//: {28}(5,900)(15,900)(15,899)(248,899){29}
//: {30}(3,898)(3,868){31}
//: {32}(5,866)(14,866)(14,867)(248,867){33}
//: {34}(3,864)(3,840){35}
//: {36}(5,838)(127,838)(127,836)(250,836){37}
//: {38}(3,836)(3,809){39}
//: {40}(5,807)(15,807)(15,803)(251,803){41}
//: {42}(3,805)(3,767){43}
//: {44}(5,765)(15,765)(15,764)(251,764){45}
//: {46}(3,763)(3,736){47}
//: {48}(5,734)(125,734)(125,733)(248,733){49}
//: {50}(3,732)(3,702){51}
//: {52}(5,700)(15,700)(15,701)(253,701){53}
//: {54}(3,698)(3,675){55}
//: {56}(5,673)(15,673)(15,669)(254,669){57}
//: {58}(3,671)(3,608){59}
//: {60}(5,606)(129,606)(129,604)(253,604){61}
//: {62}(3,604)(3,572){63}
//: {64}(5,570)(15,570)(15,572)(254,572){65}
//: {66}(3,568)(3,544){67}
//: {68}(5,542)(15,542)(15,541)(255,541){69}
//: {70}(3,540)(3,510){71}
//: {72}(5,508)(15,508)(15,509)(256,509){73}
//: {74}(3,506)(3,472){75}
//: {76}(5,470)(15,470)(15,469)(256,469){77}
//: {78}(3,468)(3,442){79}
//: {80}(5,440)(15,440)(15,437)(257,437){81}
//: {82}(3,438)(3,408){83}
//: {84}(5,406)(15,406)(15,406)(258,406){85}
//: {86}(3,404)(3,377){87}
//: {88}(5,375)(15,375)(15,374)(259,374){89}
//: {90}(3,373)(3,308){91}
//: {92}(5,306)(130,306)(130,304)(255,304){93}
//: {94}(3,304)(3,276){95}
//: {96}(5,274)(131,274)(131,272)(257,272){97}
//: {98}(3,272)(3,238){99}
//: {100}(5,236)(15,236)(15,241)(258,241){101}
//: {102}(3,234)(3,210){103}
//: {104}(5,208)(15,208)(15,209)(259,209){105}
//: {106}(3,206)(3,171){107}
//: {108}(5,169)(132,169)(132,168)(257,168){109}
//: {110}(3,167)(3,140){111}
//: {112}(5,138)(144,138)(144,137)(271,137){113}
//: {114}(3,136)(3,106){115}
//: {116}(5,104)(266,104){117}
//: {118}(3,102)(3,78){119}
//: {120}(5,76)(133,76)(133,74)(262,74){121}
//: {122}(3,74)(3,13)(87,13)(87,-15){123}
//: {124}(3,1170)(3,1199)(245,1199){125}
wire S12;    //: /sn:0 {0}(277,506)(287,506)(287,500)(517,500){1}
wire w38;    //: /sn:0 {0}(246,1177)(-75,1177)(-75,1105)(-149,1105){1}
wire w69;    //: /sn:0 {0}(946,637)(1086,637)(1086,631)(1246,631){1}
wire S24;    //: /sn:0 {0}(272,966)(547,966)(547,1023)(576,1023){1}
wire [7:0] Sa3;    //: /sn:0 {0}(#:582,1058)(892,1058)(892,766)(#:940,766){1}
wire w97;    //: /sn:0 {0}(245,1189)(73,1189)(73,1159){1}
//: {2}(75,1157)(85,1157)(85,1157)(246,1157){3}
//: {4}(73,1155)(73,1126){5}
//: {6}(75,1124)(85,1124)(85,1126)(247,1126){7}
//: {8}(73,1122)(73,1097){9}
//: {10}(75,1095)(85,1095)(85,1094)(248,1094){11}
//: {12}(73,1093)(73,1057){13}
//: {14}(75,1055)(85,1055)(85,1054)(248,1054){15}
//: {16}(73,1053)(73,1027){17}
//: {18}(75,1025)(85,1025)(85,1022)(249,1022){19}
//: {20}(73,1023)(73,993){21}
//: {22}(75,991)(85,991)(85,990)(250,990){23}
//: {24}(73,989)(73,962){25}
//: {26}(75,960)(85,960)(85,959)(251,959){27}
//: {28}(73,958)(73,894){29}
//: {30}(75,892)(85,892)(85,889)(248,889){31}
//: {32}(73,890)(73,854){33}
//: {34}(75,852)(84,852)(84,857)(248,857){35}
//: {36}(73,850)(73,823){37}
//: {38}(75,821)(85,821)(85,826)(250,826){39}
//: {40}(73,819)(73,798){41}
//: {42}(75,796)(163,796)(163,793)(251,793){43}
//: {44}(73,794)(73,754){45}
//: {46}(75,752)(85,752)(85,754)(251,754){47}
//: {48}(73,750)(73,722){49}
//: {50}(75,720)(81,720)(81,723)(248,723){51}
//: {52}(73,718)(73,694){53}
//: {54}(75,692)(85,692)(85,691)(253,691){55}
//: {56}(73,690)(73,664){57}
//: {58}(75,662)(80,662)(80,659)(254,659){59}
//: {60}(73,660)(73,595){61}
//: {62}(75,593)(85,593)(85,594)(253,594){63}
//: {64}(73,591)(73,567){65}
//: {66}(75,565)(85,565)(85,562)(254,562){67}
//: {68}(73,563)(73,539){69}
//: {70}(75,537)(85,537)(85,531)(255,531){71}
//: {72}(73,535)(73,502){73}
//: {74}(75,500)(85,500)(85,499)(256,499){75}
//: {76}(73,498)(73,463){77}
//: {78}(75,461)(165,461)(165,459)(256,459){79}
//: {80}(73,459)(73,431){81}
//: {82}(75,429)(166,429)(166,427)(257,427){83}
//: {84}(73,427)(73,398){85}
//: {86}(75,396)(85,396)(85,396)(258,396){87}
//: {88}(73,394)(73,364){89}
//: {90}(75,362)(85,362)(85,364)(259,364){91}
//: {92}(73,360)(73,300){93}
//: {94}(75,298)(84,298)(84,294)(255,294){95}
//: {96}(73,296)(73,266){97}
//: {98}(75,264)(166,264)(166,262)(257,262){99}
//: {100}(73,262)(73,236){101}
//: {102}(75,234)(85,234)(85,231)(258,231){103}
//: {104}(73,232)(73,198){105}
//: {106}(75,196)(85,196)(85,199)(259,199){107}
//: {108}(73,194)(73,163){109}
//: {110}(75,161)(174,161)(174,158)(257,158){111}
//: {112}(73,159)(73,130){113}
//: {114}(75,128)(179,128)(179,127)(271,127){115}
//: {116}(73,126)(73,96){117}
//: {118}(75,94)(266,94){119}
//: {120}(73,92)(73,70){121}
//: {122}(75,68)(85,68)(85,64)(262,64){123}
//: {124}(73,66)(73,25)(107,25)(107,-15){125}
wire [7:0] w3;    //: /sn:0 {0}(#:409,183)(878,183)(878,486)(#:940,486){1}
wire w0;    //: /sn:0 {0}(246,1162)(42,1162)(42,1159)(32,1159){1}
//: {2}(30,1157)(30,1132){3}
//: {4}(32,1130)(42,1130)(42,1131)(247,1131){5}
//: {6}(30,1128)(30,1103){7}
//: {8}(32,1101)(140,1101)(140,1099)(248,1099){9}
//: {10}(30,1099)(30,1062){11}
//: {12}(32,1060)(42,1060)(42,1059)(248,1059){13}
//: {14}(30,1058)(30,1025){15}
//: {16}(32,1023)(42,1023)(42,1027)(249,1027){17}
//: {18}(30,1021)(30,1000){19}
//: {20}(32,998)(141,998)(141,995)(250,995){21}
//: {22}(30,996)(30,966){23}
//: {24}(32,964)(42,964)(42,964)(251,964){25}
//: {26}(30,962)(30,896){27}
//: {28}(32,894)(42,894)(42,894)(248,894){29}
//: {30}(30,892)(30,864){31}
//: {32}(32,862)(41,862)(41,862)(248,862){33}
//: {34}(30,860)(30,829){35}
//: {36}(32,827)(42,827)(42,831)(250,831){37}
//: {38}(30,825)(30,803){39}
//: {40}(32,801)(141,801)(141,798)(251,798){41}
//: {42}(30,799)(30,764){43}
//: {44}(32,762)(42,762)(42,759)(251,759){45}
//: {46}(30,760)(30,732){47}
//: {48}(32,730)(38,730)(38,728)(248,728){49}
//: {50}(30,728)(30,701){51}
//: {52}(32,699)(42,699)(42,696)(253,696){53}
//: {54}(30,697)(30,668){55}
//: {56}(32,666)(143,666)(143,664)(254,664){57}
//: {58}(30,664)(30,605){59}
//: {60}(32,603)(42,603)(42,599)(253,599){61}
//: {62}(30,601)(30,569){63}
//: {64}(32,567)(42,567)(42,567)(254,567){65}
//: {66}(30,565)(30,541){67}
//: {68}(32,539)(92,539)(92,536)(255,536){69}
//: {70}(30,537)(30,504){71}
//: {72}(32,502)(42,502)(42,504)(256,504){73}
//: {74}(30,500)(30,466){75}
//: {76}(32,464)(42,464)(42,464)(256,464){77}
//: {78}(30,462)(30,436){79}
//: {80}(32,434)(144,434)(144,432)(257,432){81}
//: {82}(30,432)(30,402){83}
//: {84}(32,400)(42,400)(42,401)(258,401){85}
//: {86}(30,398)(30,373){87}
//: {88}(32,371)(145,371)(145,369)(259,369){89}
//: {90}(30,369)(30,304){91}
//: {92}(32,302)(41,302)(41,299)(255,299){93}
//: {94}(30,300)(30,271){95}
//: {96}(32,269)(144,269)(144,267)(257,267){97}
//: {98}(30,267)(30,238){99}
//: {100}(32,236)(42,236)(42,236)(258,236){101}
//: {102}(30,234)(30,208){103}
//: {104}(32,206)(145,206)(145,204)(259,204){105}
//: {106}(30,204)(30,168){107}
//: {108}(32,166)(152,166)(152,163)(257,163){109}
//: {110}(30,164)(30,137){111}
//: {112}(32,135)(53,135)(53,132)(271,132){113}
//: {114}(30,133)(30,101){115}
//: {116}(32,99)(266,99){117}
//: {118}(30,97)(30,76){119}
//: {120}(32,74)(42,74)(42,69)(262,69){121}
//: {122}(30,72)(30,19)(97,19)(97,-15){123}
//: {124}(30,1161)(30,1194)(245,1194){125}
wire w66;    //: /sn:0 {0}(946,604)(1107,604)(1107,621)(1246,621){1}
wire w64;    //: /sn:0 {0}(946,584)(1125,584)(1125,611)(1246,611){1}
wire w37;    //: /sn:0 {0}(247,1146)(-71,1146)(-71,1095)(-149,1095){1}
wire S28;    //: /sn:0 {0}(269,1101)(461,1101)(461,1063)(576,1063){1}
wire w63;    //: /sn:0 {0}(946,574)(1138,574)(1138,606)(1246,606){1}
wire w34;    //: /sn:0 {0}(249,1042)(-120,1042)(-120,1065)(-149,1065){1}
wire S26;    //: /sn:0 {0}(270,1029)(506,1029)(506,1043)(576,1043){1}
wire S18;    //: /sn:0 {0}(269,730)(484,730)(484,773)(540,773){1}
wire w76;    //: /sn:0 {0}(1246,666)(1145,666)(1145,707)(946,707){1}
wire [7:0] w43;    //: /sn:0 {0}(-421,640)(-279,640)(#:-279,467)(#:-179,467){1}
wire w21;    //: /sn:0 {0}(253,614)(-158,614)(-158,502)(-173,502){1}
wire S16;    //: /sn:0 {0}(275,666)(511,666)(511,753)(540,753){1}
wire w75;    //: /sn:0 {0}(946,697)(1138,697)(1138,661)(1246,661){1}
wire [7:0] w67;    //: /sn:0 {0}(#:-421,660)(-287,660)(-287,1080)(#:-155,1080){1}
wire S4;    //: /sn:0 {0}(403,188)(339,188)(339,206)(280,206){1}
wire S13;    //: /sn:0 {0}(276,538)(387,538)(387,510)(517,510){1}
wire w31;    //: /sn:0 {0}(946,451)(1232,451)(1232,551)(1246,551){1}
wire [7:0] w58;    //: /sn:0 {0}(#:-421,650)(-215,650)(-215,829)(#:-200,829){1}
wire S15;    //: /sn:0 {0}(274,601)(467,601)(467,530)(517,530){1}
wire w28;    //: /sn:0 {0}(250,846)(-179,846)(-179,844)(-194,844){1}
wire S9;    //: /sn:0 {0}(279,403)(472,403)(472,470)(517,470){1}
wire S8;    //: /sn:0 {0}(280,371)(488,371)(488,460)(517,460){1}
wire w24;    //: /sn:0 {0}(253,711)(-173,711)(-173,804)(-194,804){1}
wire w36;    //: /sn:0 {0}(248,1114)(-66,1114)(-66,1085)(-149,1085){1}
wire w23;    //: /sn:0 {0}(254,679)(-179,679)(-179,794)(-194,794){1}
wire w20;    //: /sn:0 {0}(254,582)(-125,582)(-125,492)(-173,492){1}
wire S17;    //: /sn:0 {0}(540,763)(497,763)(497,698)(274,698){1}
wire w1;    //: /sn:0 {0}(262,84)(-102,84)(-102,139)(-155,139){1}
wire S27;    //: /sn:0 {0}(269,1061)(453,1061)(453,1053)(576,1053){1}
wire w25;    //: /sn:0 {0}(248,743)(-162,743)(-162,814)(-194,814){1}
wire S0;    //: /sn:0 {0}(403,148)(389,148)(389,71)(283,71){1}
wire w82;    //: /sn:0 {0}(946,781)(1211,781)(1211,696)(1246,696){1}
wire w65;    //: /sn:0 {0}(946,594)(1119,594)(1119,616)(1246,616){1}
wire S5;    //: /sn:0 {0}(403,198)(353,198)(353,238)(279,238){1}
wire w74;    //: /sn:0 {0}(946,687)(1129,687)(1129,656)(1246,656){1}
wire w40;    //: /sn:0 {0}(946,461)(1223,461)(1223,556)(1246,556){1}
wire w18;    //: /sn:0 {0}(256,519)(-113,519)(-113,472)(-173,472){1}
wire w35;    //: /sn:0 {0}(248,1074)(-134,1074)(-134,1075)(-149,1075){1}
wire w8;    //: /sn:0 {0}(257,178)(-38,178)(-38,202)(-61,202)(-61,169)(-155,169){1}
wire w68;    //: /sn:0 {0}(946,614)(1088,614)(1088,626)(1246,626){1}
wire w30;    //: /sn:0 {0}(248,909)(-116,909)(-116,864)(-194,864){1}
wire w71;    //: /sn:0 {0}(946,657)(1104,657)(1104,641)(1246,641){1}
wire S21;    //: /sn:0 {0}(271,833)(470,833)(470,803)(540,803){1}
wire S30;    //: /sn:0 {0}(267,1164)(483,1164)(483,1083)(576,1083){1}
wire [7:0] w22;    //: /sn:0 {0}(#:546,788)(845,788)(845,672)(#:940,672){1}
wire w17;    //: /sn:0 {0}(256,479)(-108,479)(-108,462)(-173,462){1}
wire S20;    //: /sn:0 {0}(272,800)(458,800)(458,793)(540,793){1}
wire S14;    //: /sn:0 {0}(275,569)(445,569)(445,520)(517,520){1}
wire w84;    //: /sn:0 {0}(1246,706)(1226,706)(1226,801)(946,801){1}
wire w62;    //: /sn:0 {0}(946,564)(1146,564)(1146,601)(1246,601){1}
wire S31;    //: /sn:0 {0}(266,1196)(547,1196)(547,1093)(576,1093){1}
wire w49;    //: /sn:0 {0}(946,521)(1185,521)(1185,586)(1246,586){1}
wire w11;    //: /sn:0 {0}(258,251)(-118,251)(-118,189)(-155,189){1}
wire w44;    //: /sn:0 {0}(946,471)(1214,471)(1214,561)(1246,561){1}
wire w12;    //: /sn:0 {0}(257,282)(-127,282)(-127,199)(-155,199){1}
wire w2;    //: /sn:0 {0}(266,114)(-80,114)(-80,149)(-155,149){1}
wire w83;    //: /sn:0 {0}(1246,701)(1218,701)(1218,791)(946,791){1}
wire w77;    //: /sn:0 {0}(946,731)(1162,731)(1162,671)(1246,671){1}
wire S19;    //: /sn:0 {0}(272,761)(481,761)(481,783)(540,783){1}
wire w78;    //: /sn:0 {0}(946,741)(1170,741)(1170,676)(1246,676){1}
wire w10;    //: /sn:0 {0}(246,1172)(97,1172)(97,1174)(-51,1174){1}
//: {2}(-53,1172)(-53,1143){3}
//: {4}(-51,1141)(-41,1141)(-41,1141)(247,1141){5}
//: {6}(-53,1139)(-53,1107){7}
//: {8}(-51,1105)(-41,1105)(-41,1109)(248,1109){9}
//: {10}(-53,1103)(-53,1073){11}
//: {12}(-51,1071)(98,1071)(98,1069)(248,1069){13}
//: {14}(-53,1069)(-53,1035){15}
//: {16}(-51,1033)(-41,1033)(-41,1037)(249,1037){17}
//: {18}(-53,1031)(-53,1010){19}
//: {20}(-51,1008)(99,1008)(99,1005)(250,1005){21}
//: {22}(-53,1006)(-53,976){23}
//: {24}(-51,974)(-41,974)(-41,974)(251,974){25}
//: {26}(-53,972)(-53,907){27}
//: {28}(-51,905)(-41,905)(-41,904)(248,904){29}
//: {30}(-53,903)(-53,873){31}
//: {32}(-51,871)(-42,871)(-42,872)(248,872){33}
//: {34}(-53,869)(-53,842){35}
//: {36}(-51,840)(-41,840)(-41,841)(250,841){37}
//: {38}(-53,838)(-53,808){39}
//: {40}(-51,806)(-41,806)(-41,808)(251,808){41}
//: {42}(-53,804)(-53,773){43}
//: {44}(-51,771)(100,771)(100,769)(251,769){45}
//: {46}(-53,769)(-53,740){47}
//: {48}(-51,738)(248,738){49}
//: {50}(-53,736)(-53,704){51}
//: {52}(-51,702)(-41,702)(-41,706)(253,706){53}
//: {54}(-53,700)(-53,680){55}
//: {56}(-51,678)(-41,678)(-41,674)(254,674){57}
//: {58}(-53,676)(-53,613){59}
//: {60}(-51,611)(101,611)(101,609)(253,609){61}
//: {62}(-53,609)(-53,577){63}
//: {64}(-51,575)(-41,575)(-41,577)(254,577){65}
//: {66}(-53,573)(-53,549){67}
//: {68}(-51,547)(-41,547)(-41,546)(255,546){69}
//: {70}(-53,545)(-53,510){71}
//: {72}(-51,508)(-41,508)(-41,514)(256,514){73}
//: {74}(-53,506)(-53,475){75}
//: {76}(-51,473)(-41,473)(-41,474)(256,474){77}
//: {78}(-53,471)(-53,444){79}
//: {80}(-51,442)(-41,442)(-41,442)(257,442){81}
//: {82}(-53,440)(-53,410){83}
//: {84}(-51,408)(-41,408)(-41,411)(258,411){85}
//: {86}(-53,406)(-53,385){87}
//: {88}(-51,383)(-41,383)(-41,379)(259,379){89}
//: {90}(-53,381)(-53,310){91}
//: {92}(-51,308)(-42,308)(-42,309)(255,309){93}
//: {94}(-53,306)(-53,280){95}
//: {96}(-51,278)(-41,278)(-41,277)(257,277){97}
//: {98}(-53,276)(-53,240){99}
//: {100}(-51,238)(-41,238)(-41,246)(258,246){101}
//: {102}(-53,236)(-53,213){103}
//: {104}(-51,211)(-41,211)(-41,214)(259,214){105}
//: {106}(-53,209)(-53,182){107}
//: {108}(-51,180)(-43,180)(-43,173)(257,173){109}
//: {110}(-53,178)(-53,144){111}
//: {112}(-51,142)(271,142){113}
//: {114}(-53,140)(-53,111){115}
//: {116}(-51,109)(266,109){117}
//: {118}(-53,107)(-53,84){119}
//: {120}(-51,82)(30,82)(30,79)(262,79){121}
//: {122}(-53,80)(-53,9)(77,9)(77,-15){123}
//: {124}(-53,1176)(-53,1204)(245,1204){125}
wire w72;    //: /sn:0 {0}(946,667)(1113,667)(1113,646)(1246,646){1}
wire w13;    //: /sn:0 {0}(255,314)(-140,314)(-140,209)(-155,209){1}
wire w27;    //: /sn:0 {0}(251,813)(-146,813)(-146,834)(-194,834){1}
wire w48;    //: /sn:0 {0}(946,511)(1190,511)(1190,581)(1246,581){1}
wire [7:0] w5;    //: /sn:0 {0}(#:523,495)(#:801,495)(801,579)(#:940,579){1}
wire w33;    //: /sn:0 {0}(250,1010)(-128,1010)(-128,1055)(-149,1055){1}
wire S22;    //: /sn:0 {0}(269,864)(471,864)(471,813)(540,813){1}
wire S10;    //: /sn:0 {0}(278,434)(453,434)(453,480)(517,480){1}
wire w95;    //: /sn:0 {0}(946,647)(1094,647)(1094,636)(1246,636){1}
wire w47;    //: /sn:0 {0}(946,501)(1195,501)(1195,576)(1246,576){1}
wire S3;    //: /sn:0 {0}(403,178)(347,178)(347,165)(278,165){1}
wire w80;    //: /sn:0 {0}(946,761)(1189,761)(1189,686)(1246,686){1}
wire w29;    //: /sn:0 {0}(248,877)(-90,877)(-90,854)(-194,854){1}
wire w79;    //: /sn:0 {0}(946,751)(1179,751)(1179,681)(1246,681){1}
wire w9;    //: /sn:0 {0}(259,219)(-113,219)(-113,179)(-155,179){1}
wire [7:0] w42;    //: /sn:0 {0}(-421,630)(-326,630)(#:-326,174)(#:-161,174){1}
wire S23;    //: /sn:0 {0}(269,896)(511,896)(511,823)(540,823){1}
wire S29;    //: /sn:0 {0}(268,1133)(469,1133)(469,1073)(576,1073){1}
wire w39;    //: /sn:0 {0}(245,1209)(-108,1209)(-108,1115)(-149,1115){1}
wire w26;    //: /sn:0 {0}(251,774)(-152,774)(-152,824)(-194,824){1}
wire S11;    //: /sn:0 {0}(277,466)(442,466)(442,490)(517,490){1}
wire S2;    //: /sn:0 {0}(292,134)(366,134)(366,168)(403,168){1}
//: enddecls

  assign {w49, w48, w47, w46, w45, w44, w40, w31} = w3; //: CONCAT g4  @(941,486) /sn:0 /R:2 /w:[ 0 0 0 0 1 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w30, w29, w28, w27, w26, w25, w24, w23} = w58; //: CONCAT g8  @(-199,829) /sn:0 /R:2 /w:[ 1 1 1 1 1 1 1 1 1 ] /dr:0 /tp:0 /drp:0
  //: joint g165 (w4) @(3, 765) /w:[ 44 46 -1 43 ]
  //: joint g154 (w4) @(3, 700) /w:[ 52 54 -1 51 ]
  assign {w76, w75, w74, w73, w72, w71, w95, w69} = w22; //: CONCAT g13  @(941,672) /sn:0 /R:2 /w:[ 1 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: joint g186 (w6) @(117, 955) /w:[ 26 28 -1 25 ]
  //: joint g140 (w10) @(-53, 575) /w:[ 64 66 -1 63 ]
  _GGAND6 #(14) g37 (.I0(w6), .I1(!w97), .I2(w0), .I3(!w4), .I4(!w10), .I5(w11), .Z(S5));   //: @(269,238) /sn:0 /w:[ 103 103 101 101 101 0 1 ]
  _GGAND6 #(14) g55 (.I0(w6), .I1(!w97), .I2(w0), .I3(w4), .I4(w10), .I5(w37), .Z(S29));   //: @(258,1133) /sn:0 /w:[ 7 7 5 5 5 0 0 ]
  _GGAND6 #(14) g58 (.I0(w6), .I1(w97), .I2(!w0), .I3(!w4), .I4(w10), .I5(w26), .Z(S19));   //: @(262,761) /sn:0 /w:[ 47 47 45 45 45 0 0 ]
  //: joint g139 (w4) @(3, 570) /w:[ 64 66 -1 63 ]
  //: joint g112 (w97) @(73, 396) /w:[ 86 88 -1 85 ]
  //: joint g211 (w6) @(117, 1124) /w:[ 6 8 -1 5 ]
  //: joint g76 (w6) @(117, 123) /w:[ 114 116 -1 113 ]
  //: joint g111 (w6) @(117, 393) /w:[ 86 88 -1 85 ]
  //: joint g218 (w0) @(30, 1159) /w:[ 1 2 -1 124 ]
  //: joint g176 (w6) @(117, 852) /w:[ 34 36 -1 33 ]
  //: joint g157 (w97) @(73, 720) /w:[ 50 52 -1 49 ]
  assign w5 = {S15, S14, S13, S12, S11, S10, S9, S8}; //: CONCAT g1  @(522,495) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: joint g163 (w97) @(73, 752) /w:[ 46 48 -1 45 ]
  _GGAND6 #(14) g64 (.I0(!w6), .I1(!w97), .I2(!w0), .I3(!w4), .I4(w10), .I5(w23), .Z(S16));   //: @(265,666) /sn:0 /w:[ 59 59 57 57 57 0 0 ]
  //: IN g11 (E) @(-586,633) /sn:0 /w:[ 0 ]
  //: joint g166 (w6) @(117, 791) /w:[ 42 44 -1 41 ]
  //: joint g206 (w6) @(117, 1091) /w:[ 10 12 -1 9 ]
  //: joint g130 (w10) @(-53, 508) /w:[ 72 74 -1 71 ]
  //: joint g121 (w97) @(73, 461) /w:[ 78 80 -1 77 ]
  _GGAND6 #(14) g50 (.I0(w6), .I1(!w97), .I2(w0), .I3(!w4), .I4(w10), .I5(w28), .Z(S21));   //: @(261,833) /sn:0 /w:[ 39 39 37 37 37 0 0 ]
  //: joint g197 (w97) @(73, 1025) /w:[ 18 20 -1 17 ]
  //: joint g132 (w6) @(117, 527) /w:[ 70 72 -1 69 ]
  //: joint g113 (w0) @(30, 400) /w:[ 84 86 -1 83 ]
  //: joint g150 (w10) @(-53, 678) /w:[ 56 58 -1 55 ]
  //: joint g146 (w97) @(73, 662) /w:[ 58 60 -1 57 ]
  assign {w13, w12, w11, w9, w8, w7, w2, w1} = w42; //: CONCAT g6  @(-160,174) /sn:0 /R:2 /w:[ 1 1 1 1 1 1 1 1 1 ] /dr:0 /tp:0 /drp:0
  //: joint g208 (w0) @(30, 1101) /w:[ 8 10 -1 7 ]
  //: joint g192 (w0) @(30, 998) /w:[ 20 22 -1 19 ]
  //: joint g177 (w0) @(30, 862) /w:[ 32 34 -1 31 ]
  _GGAND6 #(14) g38 (.I0(w6), .I1(w97), .I2(w0), .I3(!w4), .I4(!w10), .I5(w13), .Z(S7));   //: @(266,301) /sn:0 /w:[ 95 95 93 93 93 0 0 ]
  //: joint g115 (w10) @(-53, 408) /w:[ 84 86 -1 83 ]
  assign {w21, w20, w19, w18, w17, w16, w15, w14} = w43; //: CONCAT g7  @(-178,467) /sn:0 /R:2 /w:[ 1 1 1 1 1 1 1 1 1 ] /dr:0 /tp:0 /drp:0
  _GGAND6 #(14) g53 (.I0(w6), .I1(w97), .I2(w0), .I3(w4), .I4(w10), .I5(w39), .Z(S31));   //: @(256,1196) /sn:0 /w:[ 0 0 125 125 125 0 0 ]
  //: joint g75 (w10) @(-53, 109) /w:[ 116 118 -1 115 ]
  //: joint g169 (w4) @(3, 807) /w:[ 40 42 -1 39 ]
  //: joint g160 (w10) @(-53, 738) /w:[ 48 50 -1 47 ]
  //: joint g135 (w10) @(-53, 547) /w:[ 68 70 -1 67 ]
  //: joint g149 (w4) @(3, 673) /w:[ 56 58 -1 55 ]
  //: joint g124 (w4) @(3, 470) /w:[ 76 78 -1 75 ]
  //: joint g207 (w97) @(73, 1095) /w:[ 10 12 -1 9 ]
  _GGAND6 #(14) g39 (.I0(!w6), .I1(w97), .I2(w0), .I3(!w4), .I4(!w10), .I5(w12), .Z(S6));   //: @(268,269) /sn:0 /w:[ 99 99 97 97 97 0 0 ]
  //: joint g68 (w0) @(30, 74) /w:[ 120 122 -1 119 ]
  //: joint g200 (w10) @(-53, 1033) /w:[ 16 18 -1 15 ]
  _GGAND6 #(14) g48 (.I0(!w6), .I1(!w97), .I2(!w0), .I3(w4), .I4(!w10), .I5(w14), .Z(S8));   //: @(270,371) /sn:0 /w:[ 91 91 89 89 89 0 0 ]
  //: joint g195 (w10) @(-53, 1008) /w:[ 20 22 -1 19 ]
  //: joint g205 (w10) @(-53, 1071) /w:[ 12 14 -1 11 ]
  //: joint g179 (w4) @(3, 866) /w:[ 32 34 -1 31 ]
  _GGAND6 #(14) g52 (.I0(!w6), .I1(w97), .I2(w0), .I3(!w4), .I4(w10), .I5(w29), .Z(S22));   //: @(259,864) /sn:0 /w:[ 35 35 33 33 33 0 0 ]
  //: joint g106 (w6) @(117, 359) /w:[ 90 92 -1 89 ]
  //: joint g107 (w0) @(30, 371) /w:[ 88 90 -1 87 ]
  //: joint g174 (w4) @(3, 838) /w:[ 36 38 -1 35 ]
  //: joint g83 (w0) @(30, 166) /w:[ 108 110 -1 107 ]
  assign w3 = {S7, S6, S5, S4, S3, S2, S1, S0}; //: CONCAT g221  @(408,183) /sn:0 /w:[ 0 1 1 0 0 0 1 0 0 ] /dr:1 /tp:0 /drp:1
  //: joint g201 (w6) @(117, 1051) /w:[ 14 16 -1 13 ]
  //: joint g100 (w10) @(-53, 278) /w:[ 96 98 -1 95 ]
  assign {w84, w83, w82, w81, w80, w79, w78, w77} = Sa3; //: CONCAT g14  @(941,766) /sn:0 /R:2 /w:[ 1 1 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: joint g202 (w97) @(73, 1055) /w:[ 14 16 -1 13 ]
  //: joint g193 (w97) @(73, 991) /w:[ 22 24 -1 21 ]
  _GGAND6 #(14) g44 (.I0(!w6), .I1(w97), .I2(w0), .I3(w4), .I4(!w10), .I5(w20), .Z(S14));   //: @(265,569) /sn:0 /w:[ 67 67 65 65 65 0 0 ]
  _GGAND6 #(14) g47 (.I0(!w6), .I1(w97), .I2(!w0), .I3(w4), .I4(!w10), .I5(w16), .Z(S10));   //: @(268,434) /sn:0 /w:[ 83 83 81 81 81 0 0 ]
  //: joint g80 (w10) @(-53, 142) /w:[ 112 114 -1 111 ]
  //: joint g94 (w4) @(3, 236) /w:[ 100 102 -1 99 ]
  //: joint g172 (w97) @(73, 821) /w:[ 38 40 -1 37 ]
  //: joint g159 (w4) @(3, 734) /w:[ 48 50 -1 47 ]
  //: joint g84 (w4) @(3, 169) /w:[ 108 110 -1 107 ]
  //: joint g105 (w10) @(-53, 308) /w:[ 92 94 -1 91 ]
  //: joint g155 (w10) @(-53, 702) /w:[ 52 54 -1 51 ]
  //: joint g141 (w6) @(117, 586) /w:[ 62 64 -1 61 ]
  _GGAND6 #(14) g41 (.I0(w6), .I1(!w97), .I2(!w0), .I3(w4), .I4(!w10), .I5(w15), .Z(S9));   //: @(269,403) /sn:0 /w:[ 87 87 85 85 85 0 0 ]
  //: joint g151 (w6) @(117, 687) /w:[ 54 56 -1 53 ]
  _GGAND6 #(14) g40 (.I0(!w6), .I1(!w97), .I2(w0), .I3(!w4), .I4(!w10), .I5(w9), .Z(S4));   //: @(270,206) /sn:0 /w:[ 107 107 105 105 105 0 1 ]
  _GGAND6 #(14) g54 (.I0(!w6), .I1(!w97), .I2(!w0), .I3(w4), .I4(w10), .I5(w32), .Z(S24));   //: @(262,966) /sn:0 /w:[ 27 27 25 25 25 0 0 ]
  //: joint g93 (w0) @(30, 236) /w:[ 100 102 -1 99 ]
  //: joint g116 (w6) @(117, 426) /w:[ 82 84 -1 81 ]
  //: joint g123 (w0) @(30, 464) /w:[ 76 78 -1 75 ]
  //: joint g167 (w97) @(73, 796) /w:[ 42 44 -1 41 ]
  //: IN g0 (C) @(94,-108) /sn:0 /R:3 /w:[ 1 ]
  _GGAND6 #(14) g46 (.I0(!w6), .I1(!w97), .I2(w0), .I3(w4), .I4(!w10), .I5(w18), .Z(S12));   //: @(267,506) /sn:0 /w:[ 75 75 73 73 73 0 0 ]
  //: joint g90 (w10) @(-53, 211) /w:[ 104 106 -1 103 ]
  //: joint g82 (w97) @(73, 161) /w:[ 110 112 -1 109 ]
  //: joint g136 (w6) @(117, 556) /w:[ 66 68 -1 65 ]
  //: joint g128 (w4) @(3, 508) /w:[ 72 74 -1 71 ]
  //: joint g190 (w10) @(-53, 974) /w:[ 24 26 -1 23 ]
  //: joint g173 (w0) @(30, 827) /w:[ 36 38 -1 35 ]
  _GGAND6 #(14) g33 (.I0(!w6), .I1(!w97), .I2(!w0), .I3(!w4), .I4(!w10), .I5(w1), .Z(S0));   //: @(273,71) /sn:0 /w:[ 123 123 121 121 121 0 1 ]
  //: joint g91 (w97) @(73, 234) /w:[ 102 104 -1 101 ]
  _GGAND6 #(14) g49 (.I0(w6), .I1(!w97), .I2(!w0), .I3(!w4), .I4(w10), .I5(w24), .Z(S17));   //: @(264,698) /sn:0 /w:[ 55 55 53 53 53 0 1 ]
  //: joint g198 (w0) @(30, 1023) /w:[ 16 18 -1 15 ]
  //: joint g137 (w97) @(73, 565) /w:[ 66 68 -1 65 ]
  _GGAND6 #(14) g61 (.I0(!w6), .I1(w97), .I2(!w0), .I3(!w4), .I4(w10), .I5(w25), .Z(S18));   //: @(259,730) /sn:0 /w:[ 51 51 49 49 49 0 0 ]
  assign Sa3 = {S31, S30, S29, S28, S27, S26, S25, S24}; //: CONCAT g3  @(581,1058) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: joint g220 (w4) @(3, 1168) /w:[ 1 2 -1 124 ]
  //: joint g158 (w0) @(30, 730) /w:[ 48 50 -1 47 ]
  _GGAND6 #(14) g34 (.I0(w6), .I1(!w97), .I2(!w0), .I3(!w4), .I4(!w10), .I5(w2), .Z(S1));   //: @(277,101) /sn:0 /w:[ 119 119 117 117 117 0 1 ]
  _GGAND6 #(14) g51 (.I0(w6), .I1(w97), .I2(w0), .I3(!w4), .I4(w10), .I5(w30), .Z(S23));   //: @(259,896) /sn:0 /w:[ 31 31 29 29 29 0 0 ]
  //: joint g86 (w6) @(117, 193) /w:[ 106 108 -1 105 ]
  //: joint g217 (w97) @(73, 1157) /w:[ 2 4 -1 1 ]
  //: joint g89 (w4) @(3, 208) /w:[ 104 106 -1 103 ]
  assign w22 = {S23, S22, S21, S20, S19, S18, S17, S16}; //: CONCAT g2  @(545,788) /sn:0 /w:[ 0 1 1 1 1 1 1 0 1 ] /dr:1 /tp:0 /drp:1
  assign {w10, w4, w0, w97, w6} = C; //: CONCAT g65  @(97,-20) /sn:0 /R:1 /w:[ 123 123 123 125 125 0 ] /dr:0 /tp:0 /drp:0
  //: joint g77 (w97) @(73, 128) /w:[ 114 116 -1 113 ]
  //: joint g110 (w10) @(-53, 383) /w:[ 88 90 -1 87 ]
  //: joint g213 (w0) @(30, 1130) /w:[ 4 6 -1 3 ]
  //: joint g156 (w6) @(117, 717) /w:[ 50 52 -1 49 ]
  //: joint g148 (w0) @(30, 666) /w:[ 56 58 -1 55 ]
  //: joint g147 (w6) @(117, 647) /w:[ 58 60 -1 57 ]
  _GGAND6 #(14) g59 (.I0(w6), .I1(!w97), .I2(!w0), .I3(w4), .I4(w10), .I5(w33), .Z(S25));   //: @(261,997) /sn:0 /w:[ 23 23 21 21 21 0 0 ]
  //: joint g203 (w0) @(30, 1060) /w:[ 12 14 -1 11 ]
  //: joint g153 (w97) @(73, 692) /w:[ 54 56 -1 53 ]
  //: joint g72 (w97) @(73, 94) /w:[ 118 120 -1 117 ]
  //: joint g161 (w6) @(117, 752) /w:[ 46 48 -1 45 ]
  //: joint g182 (w97) @(73, 892) /w:[ 30 32 -1 29 ]
  //: joint g99 (w4) @(3, 274) /w:[ 96 98 -1 95 ]
  //: joint g98 (w0) @(30, 269) /w:[ 96 98 -1 95 ]
  //: joint g196 (w6) @(117, 1020) /w:[ 18 20 -1 17 ]
  //: joint g96 (w6) @(117, 259) /w:[ 98 100 -1 97 ]
  //: joint g189 (w4) @(3, 969) /w:[ 24 26 -1 23 ]
  //: joint g183 (w0) @(30, 894) /w:[ 28 30 -1 27 ]
  //: joint g152 (w0) @(30, 699) /w:[ 52 54 -1 51 ]
  //: joint g103 (w0) @(30, 302) /w:[ 92 94 -1 91 ]
  //: joint g122 (w6) @(117, 454) /w:[ 78 80 -1 77 ]
  //: joint g87 (w97) @(73, 196) /w:[ 106 108 -1 105 ]
  //: joint g78 (w0) @(30, 135) /w:[ 112 114 -1 111 ]
  //: joint g212 (w97) @(73, 1124) /w:[ 6 8 -1 5 ]
  assign {w67, w58, w43, w42} = E; //: CONCAT g10  @(-426,645) /sn:0 /R:2 /w:[ 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: joint g129 (w0) @(30, 502) /w:[ 72 74 -1 71 ]
  //: joint g171 (w6) @(117, 823) /w:[ 38 40 -1 37 ]
  //: joint g199 (w4) @(3, 1028) /w:[ 16 18 -1 15 ]
  //: joint g102 (w97) @(73, 298) /w:[ 94 96 -1 93 ]
  //: joint g187 (w0) @(30, 964) /w:[ 24 26 -1 23 ]
  //: joint g69 (w4) @(3, 76) /w:[ 120 122 -1 119 ]
  //: joint g143 (w0) @(30, 603) /w:[ 60 62 -1 59 ]
  //: joint g119 (w4) @(3, 440) /w:[ 80 82 -1 79 ]
  _GGAND6 #(14) g57 (.I0(!w6), .I1(w97), .I2(!w0), .I3(w4), .I4(w10), .I5(w34), .Z(S26));   //: @(260,1029) /sn:0 /w:[ 19 19 17 17 17 0 0 ]
  assign {w39, w38, w37, w36, w35, w34, w33, w32} = w67; //: CONCAT g9  @(-154,1080) /sn:0 /R:2 /w:[ 1 1 1 1 1 1 1 1 1 ] /dr:0 /tp:0 /drp:0
  //: joint g71 (w6) @(117, 92) /w:[ 118 120 -1 117 ]
  //: joint g142 (w97) @(73, 593) /w:[ 62 64 -1 61 ]
  //: OUT g15 (Sa) @(1360,628) /sn:0 /w:[ 1 ]
  //: joint g162 (w0) @(30, 762) /w:[ 44 46 -1 43 ]
  //: joint g127 (w97) @(73, 500) /w:[ 74 76 -1 73 ]
  //: joint g67 (w97) @(73, 68) /w:[ 122 124 -1 121 ]
  //: joint g131 (w97) @(73, 537) /w:[ 70 72 -1 69 ]
  _GGAND6 #(14) g43 (.I0(w6), .I1(w97), .I2(w0), .I3(w4), .I4(!w10), .I5(w21), .Z(S15));   //: @(264,601) /sn:0 /w:[ 63 63 61 61 61 0 0 ]
  //: joint g104 (w4) @(3, 306) /w:[ 92 94 -1 91 ]
  //: joint g88 (w0) @(30, 206) /w:[ 104 106 -1 103 ]
  //: joint g73 (w0) @(30, 99) /w:[ 116 118 -1 115 ]
  _GGAND6 #(14) g62 (.I0(w6), .I1(w97), .I2(!w0), .I3(w4), .I4(w10), .I5(w35), .Z(S27));   //: @(259,1061) /sn:0 /w:[ 15 15 13 13 13 0 0 ]
  //: joint g145 (w10) @(-53, 611) /w:[ 60 62 -1 59 ]
  _GGAND6 #(14) g63 (.I0(!w6), .I1(!w97), .I2(w0), .I3(w4), .I4(w10), .I5(w36), .Z(S28));   //: @(259,1101) /sn:0 /w:[ 11 11 9 9 9 0 0 ]
  _GGAND6 #(14) g42 (.I0(w6), .I1(!w97), .I2(w0), .I3(w4), .I4(!w10), .I5(w19), .Z(S13));   //: @(266,538) /sn:0 /w:[ 71 71 69 69 69 0 0 ]
  //: joint g138 (w0) @(30, 567) /w:[ 64 66 -1 63 ]
  //: joint g180 (w10) @(-53, 871) /w:[ 32 34 -1 31 ]
  //: joint g188 (w97) @(73, 960) /w:[ 26 28 -1 25 ]
  //: joint g109 (w4) @(3, 375) /w:[ 88 90 -1 87 ]
  //: joint g74 (w4) @(3, 104) /w:[ 116 118 -1 115 ]
  //: joint g175 (w10) @(-53, 840) /w:[ 36 38 -1 35 ]
  _GGAND6 #(14) g56 (.I0(!w6), .I1(w97), .I2(w0), .I3(w4), .I4(w10), .I5(w38), .Z(S30));   //: @(257,1164) /sn:0 /w:[ 3 3 0 0 0 0 0 ]
  //: joint g133 (w0) @(30, 539) /w:[ 68 70 -1 67 ]
  //: joint g168 (w0) @(30, 801) /w:[ 40 42 -1 39 ]
  //: joint g181 (w6) @(117, 885) /w:[ 30 32 -1 29 ]
  _GGOR32 #(66) g5 (.I0(w31), .I1(w40), .I2(w44), .I3(w45), .I4(w46), .I5(w47), .I6(w48), .I7(w49), .I8(w60), .I9(w61), .I10(w62), .I11(w63), .I12(w64), .I13(w65), .I14(w66), .I15(w68), .I16(w69), .I17(w95), .I18(w71), .I19(w72), .I20(w73), .I21(w74), .I22(w75), .I23(w76), .I24(w77), .I25(w78), .I26(w79), .I27(w80), .I28(w81), .I29(w82), .I30(w83), .I31(w84), .Z(Sa));   //: @(1257,628) /sn:0 /w:[ 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 0 ]
  //: joint g117 (w97) @(73, 429) /w:[ 82 84 -1 81 ]
  //: joint g95 (w10) @(-53, 238) /w:[ 100 102 -1 99 ]
  //: joint g79 (w4) @(3, 138) /w:[ 112 114 -1 111 ]
  //: joint g194 (w4) @(3, 1002) /w:[ 20 22 -1 19 ]
  //: joint g215 (w10) @(-53, 1141) /w:[ 4 6 -1 3 ]
  //: joint g92 (w6) @(117, 228) /w:[ 102 104 -1 101 ]
  //: joint g85 (w10) @(-53, 180) /w:[ 108 110 -1 107 ]
  _GGAND6 #(14) g36 (.I0(w6), .I1(w97), .I2(!w0), .I3(!w4), .I4(!w10), .I5(w8), .Z(S3));   //: @(268,165) /sn:0 /w:[ 111 111 109 109 109 0 1 ]
  //: joint g216 (w6) @(117, 1151) /w:[ 2 4 -1 1 ]
  //: joint g125 (w10) @(-53, 473) /w:[ 76 78 -1 75 ]
  //: joint g144 (w4) @(3, 606) /w:[ 60 62 -1 59 ]
  //: joint g178 (w97) @(73, 852) /w:[ 34 36 -1 33 ]
  //: joint g101 (w6) @(117, 292) /w:[ 94 96 -1 93 ]
  //: joint g81 (w6) @(117, 156) /w:[ 110 112 -1 109 ]
  _GGAND6 #(14) g60 (.I0(!w6), .I1(!w97), .I2(w0), .I3(!w4), .I4(w10), .I5(w27), .Z(S20));   //: @(262,800) /sn:0 /w:[ 43 43 41 41 41 0 0 ]
  //: joint g210 (w10) @(-53, 1105) /w:[ 8 10 -1 7 ]
  //: joint g214 (w4) @(3, 1135) /w:[ 4 6 -1 3 ]
  //: joint g126 (w6) @(117, 496) /w:[ 74 76 -1 73 ]
  //: joint g70 (w10) @(-53, 82) /w:[ 120 122 -1 119 ]
  _GGAND6 #(14) g45 (.I0(w6), .I1(w97), .I2(!w0), .I3(w4), .I4(!w10), .I5(w17), .Z(S11));   //: @(267,466) /sn:0 /w:[ 79 79 77 77 77 0 0 ]
  _GGAND6 #(14) g35 (.I0(!w6), .I1(w97), .I2(!w0), .I3(!w4), .I4(!w10), .I5(w7), .Z(S2));   //: @(282,134) /sn:0 /w:[ 115 115 113 113 113 0 0 ]
  //: joint g170 (w10) @(-53, 806) /w:[ 40 42 -1 39 ]
  //: joint g185 (w10) @(-53, 905) /w:[ 28 30 -1 27 ]
  //: joint g204 (w4) @(3, 1064) /w:[ 12 14 -1 11 ]
  //: joint g120 (w10) @(-53, 442) /w:[ 80 82 -1 79 ]
  //: joint g114 (w4) @(3, 406) /w:[ 84 86 -1 83 ]
  //: joint g97 (w97) @(73, 264) /w:[ 98 100 -1 97 ]
  //: joint g66 (w6) @(117, 62) /w:[ 122 124 -1 121 ]
  //: joint g184 (w4) @(3, 900) /w:[ 28 30 -1 27 ]
  //: joint g209 (w4) @(3, 1106) /w:[ 8 10 -1 7 ]
  assign {w68, w66, w65, w64, w63, w62, w61, w60} = w5; //: CONCAT g12  @(941,579) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: joint g108 (w97) @(73, 362) /w:[ 90 92 -1 89 ]
  //: joint g164 (w10) @(-53, 771) /w:[ 44 46 -1 43 ]
  //: joint g191 (w6) @(117, 988) /w:[ 22 24 -1 21 ]
  //: joint g219 (w10) @(-53, 1174) /w:[ 1 2 -1 124 ]
  //: joint g118 (w0) @(30, 434) /w:[ 80 82 -1 79 ]
  //: joint g134 (w4) @(3, 542) /w:[ 68 70 -1 67 ]

endmodule
//: /netlistEnd

//: /netlistBegin Mux5x32
module Mux5x32(E15, C, E18, E6, E5, E1, E28, E27, E25, E16, E7, E31, E4, E0, E17, E2, E12, E29, E3, E24, E23, E9, E8, E21, E14, E13, E30, E22, E10, E19, Sa, E26, E11, E20);
//: interface  /sz:(40, 835) /bd:[ Ti0>C[4:0](19/40) Li0>E31[31:0](785/835) Li1>E30[31:0](761/835) Li2>E29[31:0](736/835) Li3>E28[31:0](712/835) Li4>E27[31:0](687/835) Li5>E26[31:0](663/835) Li6>E25[31:0](638/835) Li7>E24[31:0](613/835) Li8>E23[31:0](589/835) Li9>E22[31:0](564/835) Li10>E21[31:0](540/835) Li11>E20[31:0](515/835) Li12>E19[31:0](491/835) Li13>E18[31:0](466/835) Li14>E17[31:0](442/835) Li15>E16[31:0](417/835) Li16>E15[31:0](392/835) Li17>E14[31:0](368/835) Li18>E13[31:0](343/835) Li19>E12[31:0](319/835) Li20>E11[31:0](294/835) Li21>E10[31:0](270/835) Li22>E9[31:0](245/835) Li23>E8[31:0](221/835) Li24>E7[31:0](196/835) Li25>E6[31:0](171/835) Li26>E5[31:0](147/835) Li27>E4[31:0](122/835) Li28>E3[31:0](98/835) Li29>E2[31:0](73/835) Li30>E1[31:0](49/835) Li31>E0[31:0](24/835) Ro0<Sa[31:0](358/835) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [31:0] E12;    //: /sn:0 {0}(#:267,114)(287,114)(287,113)(302,113){1}
input [31:0] E7;    //: /sn:0 {0}(#:259,-53)(302,-53){1}
input [31:0] E20;    //: /sn:0 {0}(#:257,381)(287,381)(287,380)(302,380){1}
input [31:0] E18;    //: /sn:0 {0}(#:259,311)(287,311)(287,313)(302,313){1}
input [31:0] E29;    //: /sn:0 {0}(#:252,682)(287,682)(287,680)(302,680){1}
input [31:0] E24;    //: /sn:0 {0}(#:253,512)(287,512)(287,513)(302,513){1}
input [31:0] E10;    //: /sn:0 {0}(#:265,48)(287,48)(287,47)(302,47){1}
input [31:0] E1;    //: /sn:0 {0}(#:264,-253)(302,-253){1}
input [31:0] E19;    //: /sn:0 {0}(#:256,348)(287,348)(287,347)(302,347){1}
input [31:0] E23;    //: /sn:0 {0}(#:252,479)(287,479)(287,480)(302,480){1}
input [31:0] E21;    //: /sn:0 {0}(#:254,412)(287,412)(287,413)(302,413){1}
input [31:0] E2;    //: /sn:0 {0}(#:264,-220)(302,-220){1}
input [31:0] E30;    //: /sn:0 {0}(302,713)(268,713)(268,709)(#:261,709){1}
input [31:0] E25;    //: /sn:0 {0}(#:259,543)(287,543)(287,546)(302,546){1}
input [31:0] E0;    //: /sn:0 {0}(#:266,-285)(287,-285)(287,-286)(302,-286){1}
input [31:0] E31;    //: /sn:0 {0}(#:255,742)(287,742)(287,746)(302,746){1}
input [31:0] E16;    //: /sn:0 {0}(#:253,247)(302,247){1}
input [31:0] E14;    //: /sn:0 {0}(#:263,180)(302,180){1}
input [31:0] E28;    //: /sn:0 {0}(#:259,645)(287,645)(287,646)(302,646){1}
input [31:0] E22;    //: /sn:0 {0}(#:257,443)(287,443)(287,446)(302,446){1}
input [31:0] E13;    //: /sn:0 {0}(#:258,147)(302,147){1}
input [31:0] E8;    //: /sn:0 {0}(#:257,-20)(302,-20){1}
output [31:0] Sa;    //: /sn:0 {0}(#:1404,244)(1473,244){1}
input [31:0] E4;    //: /sn:0 {0}(#:261,-152)(277,-152)(277,-153)(302,-153){1}
input [31:0] E3;    //: /sn:0 {0}(#:258,-188)(279,-188)(279,-186)(302,-186){1}
input [4:0] C;    //: /sn:0 {0}(#:690,528)(690,525)(581,525){1}
//: {2}(579,523)(579,498){3}
//: {4}(579,494)(579,460){5}
//: {6}(581,458)(690,458)(#:690,462){7}
//: {8}(579,456)(579,434){9}
//: {10}(579,430)(579,393){11}
//: {12}(581,391)(690,391)(#:690,395){13}
//: {14}(579,389)(579,361){15}
//: {16}(579,357)(579,325){17}
//: {18}(581,323)(690,323)(#:690,328){19}
//: {20}(579,321)(579,292){21}
//: {22}(579,288)(579,262){23}
//: {24}(581,260)(690,260)(#:690,262){25}
//: {26}(579,258)(579,227){27}
//: {28}(579,223)(579,193){29}
//: {30}(581,191)(703,191)(#:703,196){31}
//: {32}(579,189)(579,160){33}
//: {34}(579,156)(579,125){35}
//: {36}(581,123)(703,123)(#:703,129){37}
//: {38}(579,121)(579,91){39}
//: {40}(579,87)(579,63){41}
//: {42}(581,61)(670,61)(670,55)(703,55)(#:703,62){43}
//: {44}(579,59)(579,23){45}
//: {46}(579,19)(579,-6){47}
//: {48}(581,-8)(703,-8)(#:703,-4){49}
//: {50}(579,-10)(579,-39){51}
//: {52}(579,-43)(579,-75){53}
//: {54}(581,-77)(703,-77)(#:703,-70){55}
//: {56}(579,-79)(579,-105){57}
//: {58}(579,-109)(579,-135){59}
//: {60}(581,-137)(642,-137)(642,-147)(703,-147)(#:703,-137){61}
//: {62}(579,-139)(579,-173){63}
//: {64}(579,-177)(579,-203){65}
//: {66}(581,-205)(703,-205)(#:703,-203){67}
//: {68}(579,-207)(579,-242){69}
//: {70}(579,-246)(579,-272){71}
//: {72}(581,-274)(703,-274)(#:703,-270){73}
//: {74}(579,-276)(579,-330){75}
//: {76}(579,-334)(#:579,-464){77}
//: {78}(577,-332)(418,-332)(#:418,-304){79}
//: {80}(577,-244)(418,-244)(#:418,-238){81}
//: {82}(577,-175)(418,-175)(#:418,-171){83}
//: {84}(577,-107)(418,-107)(#:418,-104){85}
//: {86}(577,-41)(418,-41)(#:418,-38){87}
//: {88}(577,21)(418,21)(#:418,28){89}
//: {90}(577,89)(418,89)(#:418,95){91}
//: {92}(577,158)(418,158)(#:418,162){93}
//: {94}(577,225)(422,225)(#:422,229){95}
//: {96}(577,290)(422,290)(#:422,295){97}
//: {98}(577,359)(422,359)(#:422,362){99}
//: {100}(577,432)(476,432)(476,421)(422,421)(#:422,429){101}
//: {102}(577,496)(495,496)(495,489)(422,489)(#:422,495){103}
//: {104}(579,527)(579,555){105}
//: {106}(577,557)(422,557)(#:422,561){107}
//: {108}(579,559)(579,589){109}
//: {110}(581,591)(690,591)(#:690,594){111}
//: {112}(579,593)(579,623){113}
//: {114}(577,625)(422,625)(#:422,628){115}
//: {116}(579,627)(579,656){117}
//: {118}(581,658)(690,658)(#:690,661){119}
//: {120}(579,660)(579,691){121}
//: {122}(577,693)(422,693)(#:422,695){123}
//: {124}(579,695)(579,727)(690,727)(#:690,728){125}
input [31:0] E5;    //: /sn:0 {0}(#:263,-120)(302,-120){1}
input [31:0] E15;    //: /sn:0 {0}(#:264,213)(302,213){1}
input [31:0] E27;    //: /sn:0 {0}(#:258,618)(287,618)(287,613)(302,613){1}
input [31:0] E11;    //: /sn:0 {0}(#:265,80)(302,80){1}
input [31:0] E6;    //: /sn:0 {0}(#:261,-86)(302,-86){1}
input [31:0] E26;    //: /sn:0 {0}(#:254,578)(287,578)(287,580)(302,580){1}
input [31:0] E9;    //: /sn:0 {0}(#:255,13)(274,13)(274,14)(302,14){1}
input [31:0] E17;    //: /sn:0 {0}(#:255,279)(287,279)(287,280)(302,280){1}
wire [31:0] w32;    //: /sn:0 {0}(350,746)(511,746)(511,746)(#:670,746){1}
wire [31:0] w45;    //: /sn:0 {0}(350,313)(374,313)(374,313)(#:402,313){1}
wire w96;    //: /sn:0 {0}(725,16)(985,16)(985,93)(1014,93){1}
wire w93;    //: /sn:0 {0}(725,216)(1000,216)(1000,153)(1014,153){1}
wire [31:0] w46;    //: /sn:0 {0}(350,280)(508,280)(508,280)(#:670,280){1}
wire [31:0] w60;    //: /sn:0 {0}(350,-186)(668,-186)(#:668,-185)(#:683,-185){1}
wire [31:0] w61;    //: /sn:0 {0}(350,-220)(#:398,-220){1}
wire w99;    //: /sn:0 {0}(440,-18)(1000,-18)(1000,83)(1014,83){1}
wire w141;    //: /sn:0 {0}(712,748)(1003,748)(1003,676)(1027,676){1}
wire [31:0] w56;    //: /sn:0 {0}(350,-53)(668,-53)(#:668,-52)(#:683,-52){1}
wire w153;    //: /sn:0 {0}(444,648)(953,648)(953,646)(1027,646){1}
wire w135;    //: /sn:0 {0}(444,315)(986,315)(986,360)(1027,360){1}
wire w81;    //: /sn:0 {0}(440,-151)(887,-151)(887,-171)(1014,-171){1}
wire [31:0] w38;    //: /sn:0 {0}(350,546)(512,546)(512,546)(#:670,546){1}
wire w129;    //: /sn:0 {0}(444,382)(965,382)(965,380)(1027,380){1}
wire [31:0] w51;    //: /sn:0 {0}(350,113)(373,113)(373,113)(#:398,113){1}
wire w69;    //: /sn:0 {0}(725,-250)(988,-250)(988,-201)(1014,-201){1}
wire w114;    //: /sn:0 {0}(712,348)(975,348)(975,370)(1027,370){1}
wire w120;    //: /sn:0 {0}(712,282)(999,282)(999,350)(1027,350){1}
wire [31:0] w37;    //: /sn:0 {0}(350,580)(387,580)(#:387,579)(#:402,579){1}
wire w66;    //: /sn:0 {0}(440,-284)(999,-284)(999,-211)(1014,-211){1}
wire w111;    //: /sn:0 {0}(440,48)(977,48)(977,103)(1014,103){1}
wire w159;    //: /sn:0 {0}(444,581)(963,581)(963,626)(1027,626){1}
wire [31:0] w34;    //: /sn:0 {0}(350,680)(655,680)(#:655,679)(#:670,679){1}
wire [31:0] w63;    //: /sn:0 {0}(350,-286)(#:398,-286){1}
wire w75;    //: /sn:0 {0}(440,-218)(978,-218)(978,-191)(1014,-191){1}
wire [31:0] w43;    //: /sn:0 {0}(350,380)(374,380)(374,380)(#:402,380){1}
wire w87;    //: /sn:0 {0}(440,-84)(970,-84)(970,-151)(1014,-151){1}
wire w102;    //: /sn:0 {0}(725,149)(924,149)(924,133)(1014,133){1}
wire [7:0] w119;    //: /sn:0 {0}(#:1398,249)(1048,249)(1048,375)(#:1033,375){1}
wire [31:0] w54;    //: /sn:0 {0}(#:683,14)(350,14){1}
wire w90;    //: /sn:0 {0}(725,82)(960,82)(960,113)(1014,113){1}
wire [31:0] w58;    //: /sn:0 {0}(350,-119)(#:683,-119){1}
wire w156;    //: /sn:0 {0}(444,715)(982,715)(982,666)(1027,666){1}
wire [31:0] w36;    //: /sn:0 {0}(350,613)(655,613)(#:655,612)(#:670,612){1}
wire [31:0] w41;    //: /sn:0 {0}(350,446)(387,446)(#:387,447)(#:402,447){1}
wire w132;    //: /sn:0 {0}(444,449)(986,449)(986,400)(1027,400){1}
wire w108;    //: /sn:0 {0}(440,182)(953,182)(953,143)(1014,143){1}
wire w126;    //: /sn:0 {0}(712,415)(973,415)(973,390)(1027,390){1}
wire [7:0] w74;    //: /sn:0 {0}(1398,239)(1041,239)(1041,118)(#:1020,118){1}
wire [31:0] w35;    //: /sn:0 {0}(350,646)(378,646)(378,646)(#:402,646){1}
wire [31:0] w40;    //: /sn:0 {0}(350,480)(507,480)(507,480)(#:670,480){1}
wire [7:0] w71;    //: /sn:0 {0}(1398,229)(1258,229)(1258,-176)(#:1020,-176){1}
wire w144;    //: /sn:0 {0}(712,548)(983,548)(983,616)(1027,616){1}
wire [7:0] w146;    //: /sn:0 {0}(#:1033,641)(1187,641)(1187,259)(#:1398,259){1}
wire [31:0] w53;    //: /sn:0 {0}(350,47)(383,47)(#:383,46)(#:398,46){1}
wire w84;    //: /sn:0 {0}(725,-50)(998,-50)(998,-141)(1014,-141){1}
wire w117;    //: /sn:0 {0}(712,482)(1007,482)(1007,410)(1027,410){1}
wire [31:0] w59;    //: /sn:0 {0}(350,-153)(#:398,-153){1}
wire w123;    //: /sn:0 {0}(444,249)(1012,249)(1012,340)(1027,340){1}
wire [31:0] w62;    //: /sn:0 {0}(350,-253)(668,-253)(#:668,-252)(#:683,-252){1}
wire [31:0] w44;    //: /sn:0 {0}(350,347)(655,347)(#:655,346)(#:670,346){1}
wire [31:0] w49;    //: /sn:0 {0}(350,180)(373,180)(373,180)(#:398,180){1}
wire [31:0] w57;    //: /sn:0 {0}(350,-86)(#:398,-86){1}
wire w150;    //: /sn:0 {0}(712,681)(959,681)(959,656)(1027,656){1}
wire w105;    //: /sn:0 {0}(440,115)(956,115)(956,123)(1014,123){1}
wire w78;    //: /sn:0 {0}(725,-117)(910,-117)(910,-161)(1014,-161){1}
wire w72;    //: /sn:0 {0}(725,-183)(1002,-183)(1002,-181)(1014,-181){1}
wire w138;    //: /sn:0 {0}(712,614)(955,614)(955,636)(1027,636){1}
wire [31:0] w52;    //: /sn:0 {0}(350,80)(516,80)(516,80)(#:683,80){1}
wire [31:0] w33;    //: /sn:0 {0}(350,713)(378,713)(378,713)(#:402,713){1}
wire [31:0] w48;    //: /sn:0 {0}(350,213)(668,213)(#:668,214)(#:683,214){1}
wire [31:0] w47;    //: /sn:0 {0}(350,247)(374,247)(374,247)(#:402,247){1}
wire w147;    //: /sn:0 {0}(444,515)(1009,515)(1009,606)(1027,606){1}
wire [31:0] w42;    //: /sn:0 {0}(350,413)(507,413)(507,413)(#:670,413){1}
wire [31:0] w50;    //: /sn:0 {0}(350,147)(516,147)(516,147)(#:683,147){1}
wire [31:0] w39;    //: /sn:0 {0}(350,513)(378,513)(378,513)(#:402,513){1}
wire [31:0] w55;    //: /sn:0 {0}(350,-20)(373,-20)(373,-20)(#:398,-20){1}
//: enddecls

  //: joint g61 (C) @(579, 61) /w:[ 42 44 -1 41 ]
  Mux5 g8 (.C(C), .E(w56), .Sa(w84));   //: @(684, -69) /sz:(40, 40) /sn:0 /p:[ Ti0>55 Li0>1 Ro0<0 ]
  Mux5 g4 (.C(C), .E(w60), .Sa(w72));   //: @(684, -202) /sz:(40, 40) /sn:0 /p:[ Ti0>67 Li0>1 Ro0<0 ]
  //: IN g86 (E15) @(262,213) /sn:0 /w:[ 0 ]
  //: joint g58 (C) @(579, -137) /w:[ 60 62 -1 59 ]
  //: joint g55 (C) @(579, -332) /w:[ -1 76 78 75 ]
  //: joint g51 (C) @(579, -41) /w:[ -1 52 86 51 ]
  //: IN g37 (C) @(579,-466) /sn:0 /R:3 /w:[ 77 ]
  assign w74 = {w93, w108, w102, w105, w90, w111, w96, w99}; //: CONCAT g34  @(1019,118) /sn:0 /w:[ 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign w71 = {w84, w87, w78, w81, w72, w75, w69, w66}; //: CONCAT g3  @(1019,-176) /sn:0 /w:[ 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  Mux5 g13 (.C(C), .E(w55), .Sa(w99));   //: @(399, -37) /sz:(40, 40) /sn:0 /p:[ Ti0>87 Li0>1 Ro0<0 ]
  //: IN g89 (E18) @(257,311) /sn:0 /w:[ 0 ]
  //: IN g77 (E6) @(259,-86) /sn:0 /w:[ 0 ]
  //: IN g76 (E5) @(261,-120) /sn:0 /w:[ 0 ]
  //: joint g65 (C) @(579, 323) /w:[ 18 20 -1 17 ]
  Mux5 g2 (.C(C), .E(w62), .Sa(w69));   //: @(684, -269) /sz:(40, 40) /sn:0 /p:[ Ti0>73 Li0>1 Ro0<0 ]
  //: joint g59 (C) @(579, -77) /w:[ 54 56 -1 53 ]
  //: IN g72 (E1) @(262,-253) /sn:0 /w:[ 0 ]
  Mux5 g1 (.C(C), .E(w63), .Sa(w66));   //: @(399, -303) /sz:(40, 40) /sn:0 /p:[ Ti0>79 Li0>1 Ro0<0 ]
  //: IN g99 (E28) @(257,645) /sn:0 /w:[ 0 ]
  //: IN g98 (E27) @(256,618) /sn:0 /w:[ 0 ]
  //: joint g64 (C) @(579, 260) /w:[ 24 26 -1 23 ]
  //: IN g96 (E25) @(257,543) /sn:0 /w:[ 0 ]
  Mux5 g16 (.C(C), .E(w49), .Sa(w108));   //: @(399, 163) /sz:(40, 40) /sn:0 /p:[ Ti0>93 Li0>1 Ro0<0 ]
  Mux5 g11 (.C(C), .E(w48), .Sa(w93));   //: @(684, 197) /sz:(40, 40) /sn:0 /p:[ Ti0>31 Li0>1 Ro0<0 ]
  //: IN g87 (E16) @(251,247) /sn:0 /w:[ 0 ]
  //: IN g78 (E7) @(257,-53) /sn:0 /w:[ 0 ]
  //: joint g50 (C) @(579, 21) /w:[ -1 46 88 45 ]
  Mux5 g28 (.C(C), .E(w38), .Sa(w144));   //: @(671, 529) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Li0>1 Ro0<0 ]
  Mux5 g10 (.C(C), .E(w52), .Sa(w90));   //: @(684, 63) /sz:(40, 40) /sn:0 /p:[ Ti0>43 Li0>1 Ro0<0 ]
  Mux5 g32 (.C(C), .E(w33), .Sa(w156));   //: @(403, 696) /sz:(40, 40) /sn:0 /p:[ Ti0>123 Li0>1 Ro0<0 ]
  Mux5 g27 (.C(C), .E(w32), .Sa(w141));   //: @(671, 729) /sz:(40, 40) /sn:0 /p:[ Ti0>125 Li0>1 Ro0<0 ]
  Mux5 g19 (.C(C), .E(w40), .Sa(w117));   //: @(671, 463) /sz:(40, 40) /sn:0 /p:[ Ti0>7 Li0>1 Ro0<0 ]
  //: IN g102 (E31) @(253,742) /sn:0 /w:[ 0 ]
  assign Sa = {w146, w119, w74, w71}; //: CONCAT g69  @(1403,244) /sn:0 /anc:1 /w:[ 0 1 0 0 0 ] /dr:1 /tp:0 /drp:1
  //: joint g38 (C) @(579, 693) /w:[ -1 121 122 124 ]
  Mux5 g6 (.C(C), .E(w58), .Sa(w78));   //: @(684, -136) /sz:(40, 40) /sn:0 /p:[ Ti0>61 Li0>1 Ro0<0 ]
  //: IN g75 (E4) @(259,-152) /sn:0 /w:[ 0 ]
  //: joint g57 (C) @(579, -205) /w:[ 66 68 -1 65 ]
  //: joint g53 (C) @(579, -175) /w:[ -1 64 82 63 ]
  Mux5 g9 (.C(C), .E(w57), .Sa(w87));   //: @(399, -103) /sz:(40, 40) /sn:0 /p:[ Ti0>85 Li0>1 Ro0<0 ]
  Mux5 g7 (.C(C), .E(w59), .Sa(w81));   //: @(399, -170) /sz:(40, 40) /sn:0 /p:[ Ti0>83 Li0>1 Ro0<0 ]
  //: IN g71 (E0) @(264,-285) /sn:0 /w:[ 0 ]
  Mux5 g31 (.C(C), .E(w35), .Sa(w153));   //: @(403, 629) /sz:(40, 40) /sn:0 /p:[ Ti0>115 Li0>1 Ro0<0 ]
  Mux5 g20 (.C(C), .E(w46), .Sa(w120));   //: @(671, 263) /sz:(40, 40) /sn:0 /p:[ Ti0>25 Li0>1 Ro0<0 ]
  Mux5 g15 (.C(C), .E(w51), .Sa(w105));   //: @(399, 96) /sz:(40, 40) /sn:0 /p:[ Ti0>91 Li0>1 Ro0<0 ]
  //: joint g68 (C) @(579, 525) /w:[ 1 2 -1 104 ]
  //: joint g67 (C) @(579, 458) /w:[ 6 8 -1 5 ]
  //: joint g39 (C) @(579, 658) /w:[ 118 117 -1 120 ]
  //: joint g48 (C) @(579, 158) /w:[ -1 34 92 33 ]
  //: joint g43 (C) @(579, 496) /w:[ -1 4 102 3 ]
  //: IN g88 (E17) @(253,279) /sn:0 /w:[ 0 ]
  //: IN g73 (E2) @(262,-220) /sn:0 /w:[ 0 ]
  //: joint g62 (C) @(579, 123) /w:[ 36 38 -1 35 ]
  Mux5 g29 (.C(C), .E(w39), .Sa(w147));   //: @(403, 496) /sz:(40, 40) /sn:0 /p:[ Ti0>103 Li0>1 Ro0<0 ]
  Mux5 g25 (.C(C), .E(w45), .Sa(w135));   //: @(403, 296) /sz:(40, 40) /sn:0 /p:[ Ti0>97 Li0>1 Ro0<0 ]
  Mux5 g17 (.C(C), .E(w53), .Sa(w111));   //: @(399, 29) /sz:(40, 40) /sn:0 /p:[ Ti0>89 Li0>1 Ro0<0 ]
  //: joint g63 (C) @(579, 191) /w:[ 30 32 -1 29 ]
  //: joint g52 (C) @(579, -107) /w:[ -1 58 84 57 ]
  //: joint g42 (C) @(579, 557) /w:[ -1 105 106 108 ]
  //: IN g83 (E12) @(265,114) /sn:0 /w:[ 0 ]
  //: IN g100 (E29) @(250,682) /sn:0 /w:[ 0 ]
  //: IN g74 (E3) @(256,-188) /sn:0 /w:[ 0 ]
  //: joint g56 (C) @(579, -274) /w:[ 72 74 -1 71 ]
  Mux5 g14 (.C(C), .E(w50), .Sa(w102));   //: @(684, 130) /sz:(40, 40) /sn:0 /p:[ Ti0>37 Li0>1 Ro0<0 ]
  Mux5 g5 (.C(C), .E(w61), .Sa(w75));   //: @(399, -237) /sz:(40, 40) /sn:0 /p:[ Ti0>81 Li0>1 Ro0<0 ]
  //: IN g95 (E24) @(251,512) /sn:0 /w:[ 0 ]
  //: IN g94 (E23) @(250,479) /sn:0 /w:[ 0 ]
  //: IN g80 (E9) @(253,13) /sn:0 /w:[ 0 ]
  //: IN g79 (E8) @(255,-20) /sn:0 /w:[ 0 ]
  //: joint g47 (C) @(579, 225) /w:[ -1 28 94 27 ]
  //: joint g44 (C) @(579, 432) /w:[ -1 10 100 9 ]
  //: IN g92 (E21) @(252,412) /sn:0 /w:[ 0 ]
  //: IN g85 (E14) @(261,180) /sn:0 /w:[ 0 ]
  //: IN g84 (E13) @(256,147) /sn:0 /w:[ 0 ]
  assign w146 = {w141, w156, w150, w153, w138, w159, w144, w147}; //: CONCAT g36  @(1032,641) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  Mux5 g24 (.C(C), .E(w41), .Sa(w132));   //: @(403, 430) /sz:(40, 40) /sn:0 /p:[ Ti0>101 Li0>1 Ro0<0 ]
  Mux5 g21 (.C(C), .E(w47), .Sa(w123));   //: @(403, 230) /sz:(40, 40) /sn:0 /p:[ Ti0>95 Li0>1 Ro0<0 ]
  //: joint g41 (C) @(579, 625) /w:[ -1 113 114 116 ]
  Mux5 g23 (.C(C), .E(w43), .Sa(w129));   //: @(403, 363) /sz:(40, 40) /sn:0 /p:[ Ti0>99 Li0>1 Ro0<0 ]
  //: IN g101 (E30) @(259,709) /sn:0 /w:[ 1 ]
  //: IN g93 (E22) @(255,443) /sn:0 /w:[ 0 ]
  //: IN g81 (E10) @(263,48) /sn:0 /w:[ 0 ]
  //: joint g60 (C) @(579, -8) /w:[ 48 50 -1 47 ]
  //: joint g54 (C) @(579, -244) /w:[ -1 70 80 69 ]
  //: joint g40 (C) @(579, 591) /w:[ 110 109 -1 112 ]
  //: IN g90 (E19) @(254,348) /sn:0 /w:[ 0 ]
  //: OUT g70 (Sa) @(1470,244) /sn:0 /w:[ 1 ]
  //: joint g46 (C) @(579, 290) /w:[ -1 22 96 21 ]
  //: joint g45 (C) @(579, 359) /w:[ -1 16 98 15 ]
  assign w119 = {w117, w132, w126, w129, w114, w135, w120, w123}; //: CONCAT g35  @(1032,375) /sn:0 /w:[ 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  Mux5 g26 (.C(C), .E(w36), .Sa(w138));   //: @(671, 595) /sz:(40, 40) /sn:0 /p:[ Ti0>111 Li0>1 Ro0<0 ]
  Mux5 g22 (.C(C), .E(w42), .Sa(w126));   //: @(671, 396) /sz:(40, 40) /sn:0 /p:[ Ti0>13 Li0>1 Ro0<0 ]
  Mux5cableado g0 (.E0(E0), .E1(E1), .E2(E2), .E3(E3), .E4(E4), .E5(E5), .E6(E6), .E7(E7), .E8(E8), .E9(E9), .E10(E10), .E11(E11), .E12(E12), .E13(E13), .E14(E14), .E15(E15), .E16(E16), .E17(E17), .E18(E18), .E19(E19), .E20(E20), .E21(E21), .E22(E22), .E23(E23), .E24(E24), .E25(E25), .E26(E26), .E27(E27), .E28(E28), .E29(E29), .E30(E30), .E31(E31), .S0(w63), .S1(w62), .S2(w61), .S3(w60), .S4(w59), .S5(w58), .S6(w57), .S7(w56), .S8(w55), .S9(w54), .S10(w53), .S11(w52), .S12(w51), .S13(w50), .S14(w49), .S15(w48), .S16(w47), .S17(w46), .S18(w45), .S19(w44), .S20(w43), .S21(w42), .S22(w41), .S23(w40), .S24(w39), .S25(w38), .S26(w37), .S27(w36), .S28(w35), .S29(w34), .S30(w33), .S31(w32));   //: @(303, -319) /sz:(46, 1099) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>1 Li5>1 Li6>1 Li7>1 Li8>1 Li9>1 Li10>1 Li11>1 Li12>1 Li13>1 Li14>1 Li15>1 Li16>1 Li17>1 Li18>1 Li19>1 Li20>1 Li21>1 Li22>1 Li23>1 Li24>1 Li25>1 Li26>1 Li27>1 Li28>1 Li29>1 Li30>0 Li31>1 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<0 Ro6<0 Ro7<0 Ro8<0 Ro9<1 Ro10<0 Ro11<0 Ro12<0 Ro13<0 Ro14<0 Ro15<0 Ro16<0 Ro17<0 Ro18<0 Ro19<0 Ro20<0 Ro21<0 Ro22<0 Ro23<0 Ro24<0 Ro25<0 Ro26<0 Ro27<0 Ro28<0 Ro29<0 Ro30<0 Ro31<0 ]
  //: IN g97 (E26) @(252,578) /sn:0 /w:[ 0 ]
  //: IN g82 (E11) @(263,80) /sn:0 /w:[ 0 ]
  //: joint g66 (C) @(579, 391) /w:[ 12 14 -1 11 ]
  Mux5 g18 (.C(C), .E(w44), .Sa(w114));   //: @(671, 329) /sz:(40, 40) /sn:0 /p:[ Ti0>19 Li0>1 Ro0<0 ]
  Mux5 g12 (.C(C), .E(w54), .Sa(w96));   //: @(684, -3) /sz:(40, 40) /sn:0 /p:[ Ti0>49 Li0>0 Ro0<0 ]
  //: IN g91 (E20) @(255,381) /sn:0 /w:[ 0 ]
  Mux5 g33 (.C(C), .E(w37), .Sa(w159));   //: @(403, 562) /sz:(40, 40) /sn:0 /p:[ Ti0>107 Li0>1 Ro0<0 ]
  Mux5 g30 (.C(C), .E(w34), .Sa(w150));   //: @(671, 662) /sz:(40, 40) /sn:0 /p:[ Ti0>119 Li0>1 Ro0<0 ]
  //: joint g49 (C) @(579, 89) /w:[ -1 40 90 39 ]

endmodule
//: /netlistEnd

//: /netlistBegin Decodificador5
module Decodificador5(S3, S7, S12, S0, S10, S27, S18, S5, S6, S19, S30, S16, S24, S28, S13, S20, S22, C, S25, S2, S1, S15, S9, S26, S31, S8, S14, S4, S23, S21, S11, S17, S29);
//: interface  /sz:(40, 957) /bd:[ Li0>C[4:0](447/957) Ro0<S31(928/957) Ro1<S30(899/957) Ro2<S29(870/957) Ro3<S28(841/957) Ro4<S27(812/957) Ro5<S26(783/957) Ro6<S25(754/957) Ro7<S24(725/957) Ro8<S23(696/957) Ro9<S22(667/957) Ro10<S21(638/957) Ro11<S20(609/957) Ro12<S19(580/957) Ro13<S18(551/957) Ro14<S17(522/957) Ro15<S16(493/957) Ro16<S15(464/957) Ro17<S14(435/957) Ro18<S13(406/957) Ro19<S12(377/957) Ro20<S11(348/957) Ro21<S10(319/957) Ro22<S9(290/957) Ro23<S8(261/957) Ro24<S7(232/957) Ro25<S6(203/957) Ro26<S5(174/957) Ro27<S4(145/957) Ro28<S3(116/957) Ro29<S2(87/957) Ro30<S1(58/957) Ro31<S0(29/957) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output S1;    //: /sn:0 {0}(277,101)(326,101)(326,104)(345,104){1}
output S25;    //: /sn:0 {0}(271,998)(348,998)(348,1006)(362,1006){1}
output S7;    //: /sn:0 {0}(277,301)(329,301)(329,302)(343,302){1}
output S6;    //: /sn:0 {0}(278,269)(329,269)(329,272)(343,272){1}
output S12;    //: /sn:0 {0}(277,506)(382,506)(382,488)(396,488){1}
output S24;    //: /sn:0 {0}(272,966)(347,966)(347,981)(361,981){1}
output S28;    //: /sn:0 {0}(269,1101)(367,1101)(367,1088)(381,1088){1}
output S18;    //: /sn:0 {0}(273,729)(375,729)(375,737)(389,737){1}
output S26;    //: /sn:0 {0}(270,1029)(354,1029)(354,1044)(368,1044){1}
output S16;    //: /sn:0 {0}(275,666)(368,666)(368,674)(382,674){1}
output S4;    //: /sn:0 {0}(339,207)(307,207)(307,206)(280,206){1}
output S13;    //: /sn:0 {0}(276,538)(371,538)(371,530)(385,530){1}
output S15;    //: /sn:0 {0}(407,574)(346,574)(346,601)(274,601){1}
output S8;    //: /sn:0 {0}(280,371)(343,371)(343,383)(357,383){1}
output S9;    //: /sn:0 {0}(279,403)(344,403)(344,408)(358,408){1}
output S17;    //: /sn:0 {0}(274,698)(369,698)(369,699)(383,699){1}
output S27;    //: /sn:0 {0}(269,1061)(358,1061)(358,1067)(372,1067){1}
output S0;    //: /sn:0 {0}(283,71)(328,71)(328,74)(339,74){1}
output S5;    //: /sn:0 {0}(279,238)(328,238)(328,240)(342,240){1}
output S21;    //: /sn:0 {0}(271,833)(346,833)(346,827)(360,827){1}
output S20;    //: /sn:0 {0}(272,801)(345,801)(345,802)(359,802){1}
output S30;    //: /sn:0 {0}(267,1164)(374,1164)(374,1151)(388,1151){1}
output S14;    //: /sn:0 {0}(403,551)(290,551)(290,569)(275,569){1}
output S31;    //: /sn:0 {0}(266,1196)(339,1196)(339,1211)(353,1211){1}
input [4:0] C;    //: /sn:0 {0}(#:97,-21)(97,-89)(94,-89)(#:94,-106){1}
output S19;    //: /sn:0 {0}(272,761)(379,761)(379,760)(393,760){1}
output S10;    //: /sn:0 {0}(278,434)(350,434)(350,446)(364,446){1}
output S22;    //: /sn:0 {0}(270,864)(352,864)(352,865)(366,865){1}
output S3;    //: /sn:0 {0}(280,166)(349,166){1}
output S23;    //: /sn:0 {0}(269,896)(356,896)(356,888)(370,888){1}
output S29;    //: /sn:0 {0}(268,1133)(368,1133)(368,1113)(382,1113){1}
output S2;    //: /sn:0 {0}(343,140)(291,140)(291,134)(281,134){1}
output S11;    //: /sn:0 {0}(277,466)(354,466)(354,469)(368,469){1}
wire w6;    //: /sn:0 {0}(245,1186)(117,1186)(117,1153){1}
//: {2}(119,1151)(129,1151)(129,1154)(246,1154){3}
//: {4}(117,1149)(117,1126){5}
//: {6}(119,1124)(129,1124)(129,1123)(247,1123){7}
//: {8}(117,1122)(117,1093){9}
//: {10}(119,1091)(248,1091){11}
//: {12}(117,1089)(117,1053){13}
//: {14}(119,1051)(248,1051){15}
//: {16}(117,1049)(117,1022){17}
//: {18}(119,1020)(129,1020)(129,1019)(249,1019){19}
//: {20}(117,1018)(117,990){21}
//: {22}(119,988)(250,988){23}
//: {24}(117,986)(117,957){25}
//: {26}(119,955)(129,955)(129,956)(251,956){27}
//: {28}(117,953)(117,887){29}
//: {30}(119,885)(129,885)(129,886)(248,886){31}
//: {32}(117,883)(117,854){33}
//: {34}(119,852)(129,852)(129,854)(249,854){35}
//: {36}(117,850)(117,825){37}
//: {38}(119,823)(250,823){39}
//: {40}(117,821)(117,793){41}
//: {42}(119,791)(251,791){43}
//: {44}(117,789)(117,754){45}
//: {46}(119,752)(129,752)(129,751)(251,751){47}
//: {48}(117,750)(117,719){49}
//: {50}(119,717)(129,717)(129,719)(252,719){51}
//: {52}(117,715)(117,689){53}
//: {54}(119,687)(129,687)(129,688)(253,688){55}
//: {56}(117,685)(117,649){57}
//: {58}(119,647)(129,647)(129,656)(254,656){59}
//: {60}(117,645)(117,588){61}
//: {62}(119,586)(129,586)(129,591)(253,591){63}
//: {64}(117,584)(117,558){65}
//: {66}(119,556)(129,556)(129,559)(254,559){67}
//: {68}(117,554)(117,529){69}
//: {70}(119,527)(129,527)(129,528)(255,528){71}
//: {72}(117,525)(117,498){73}
//: {74}(119,496)(256,496){75}
//: {76}(117,494)(117,456){77}
//: {78}(119,454)(129,454)(129,456)(256,456){79}
//: {80}(117,452)(117,428){81}
//: {82}(119,426)(129,426)(129,424)(257,424){83}
//: {84}(117,424)(117,395){85}
//: {86}(119,393)(258,393){87}
//: {88}(117,391)(117,361){89}
//: {90}(119,359)(129,359)(129,361)(259,361){91}
//: {92}(117,357)(117,294){93}
//: {94}(119,292)(129,292)(129,291)(256,291){95}
//: {96}(117,290)(117,261){97}
//: {98}(119,259)(257,259){99}
//: {100}(117,257)(117,230){101}
//: {102}(119,228)(258,228){103}
//: {104}(117,226)(117,195){105}
//: {106}(119,193)(129,193)(129,196)(259,196){107}
//: {108}(117,191)(117,158){109}
//: {110}(119,156)(259,156){111}
//: {112}(117,154)(117,125){113}
//: {114}(119,123)(129,123)(129,124)(260,124){115}
//: {116}(117,121)(117,94){117}
//: {118}(119,92)(129,92)(129,91)(256,91){119}
//: {120}(117,90)(117,64){121}
//: {122}(119,62)(129,62)(129,61)(262,61){123}
//: {124}(117,60)(117,-15){125}
wire w4;    //: /sn:0 {0}(246,1169)(15,1169)(15,1168)(5,1168){1}
//: {2}(3,1166)(3,1137){3}
//: {4}(5,1135)(15,1135)(15,1138)(247,1138){5}
//: {6}(3,1133)(3,1108){7}
//: {8}(5,1106)(248,1106){9}
//: {10}(3,1104)(3,1066){11}
//: {12}(5,1064)(15,1064)(15,1066)(248,1066){13}
//: {14}(3,1062)(3,1030){15}
//: {16}(5,1028)(15,1028)(15,1034)(249,1034){17}
//: {18}(3,1026)(3,1004){19}
//: {20}(5,1002)(15,1002)(15,1003)(250,1003){21}
//: {22}(3,1000)(3,971){23}
//: {24}(5,969)(15,969)(15,971)(251,971){25}
//: {26}(3,967)(3,902){27}
//: {28}(5,900)(15,900)(15,901)(248,901){29}
//: {30}(3,898)(3,868){31}
//: {32}(5,866)(15,866)(15,869)(249,869){33}
//: {34}(3,864)(3,840){35}
//: {36}(5,838)(250,838){37}
//: {38}(3,836)(3,809){39}
//: {40}(5,807)(15,807)(15,806)(251,806){41}
//: {42}(3,805)(3,767){43}
//: {44}(5,765)(15,765)(15,766)(251,766){45}
//: {46}(3,763)(3,736){47}
//: {48}(5,734)(252,734){49}
//: {50}(3,732)(3,702){51}
//: {52}(5,700)(15,700)(15,703)(253,703){53}
//: {54}(3,698)(3,675){55}
//: {56}(5,673)(15,673)(15,671)(254,671){57}
//: {58}(3,671)(3,608){59}
//: {60}(5,606)(253,606){61}
//: {62}(3,604)(3,572){63}
//: {64}(5,570)(15,570)(15,574)(254,574){65}
//: {66}(3,568)(3,544){67}
//: {68}(5,542)(15,542)(15,543)(255,543){69}
//: {70}(3,540)(3,510){71}
//: {72}(5,508)(15,508)(15,511)(256,511){73}
//: {74}(3,506)(3,472){75}
//: {76}(5,470)(15,470)(15,471)(256,471){77}
//: {78}(3,468)(3,442){79}
//: {80}(5,440)(15,440)(15,439)(257,439){81}
//: {82}(3,438)(3,408){83}
//: {84}(5,406)(15,406)(15,408)(258,408){85}
//: {86}(3,404)(3,377){87}
//: {88}(5,375)(15,375)(15,376)(259,376){89}
//: {90}(3,373)(3,308){91}
//: {92}(5,306)(256,306){93}
//: {94}(3,304)(3,276){95}
//: {96}(5,274)(257,274){97}
//: {98}(3,272)(3,238){99}
//: {100}(5,236)(15,236)(15,243)(258,243){101}
//: {102}(3,234)(3,210){103}
//: {104}(5,208)(15,208)(15,211)(259,211){105}
//: {106}(3,206)(3,171){107}
//: {108}(5,169)(15,169)(15,171)(259,171){109}
//: {110}(3,167)(3,140){111}
//: {112}(5,138)(15,138)(15,139)(260,139){113}
//: {114}(3,136)(3,106){115}
//: {116}(5,104)(15,104)(15,106)(256,106){117}
//: {118}(3,102)(3,78){119}
//: {120}(5,76)(262,76){121}
//: {122}(3,74)(3,13)(87,13)(87,-15){123}
//: {124}(3,1170)(3,1201)(245,1201){125}
wire w0;    //: /sn:0 {0}(246,1164)(42,1164)(42,1159)(32,1159){1}
//: {2}(30,1157)(30,1132){3}
//: {4}(32,1130)(42,1130)(42,1133)(247,1133){5}
//: {6}(30,1128)(30,1103){7}
//: {8}(32,1101)(248,1101){9}
//: {10}(30,1099)(30,1062){11}
//: {12}(32,1060)(42,1060)(42,1061)(248,1061){13}
//: {14}(30,1058)(30,1025){15}
//: {16}(32,1023)(42,1023)(42,1029)(249,1029){17}
//: {18}(30,1021)(30,1000){19}
//: {20}(32,998)(250,998){21}
//: {22}(30,996)(30,966){23}
//: {24}(32,964)(42,964)(42,966)(251,966){25}
//: {26}(30,962)(30,896){27}
//: {28}(32,894)(42,894)(42,896)(248,896){29}
//: {30}(30,892)(30,864){31}
//: {32}(32,862)(42,862)(42,864)(249,864){33}
//: {34}(30,860)(30,829){35}
//: {36}(32,827)(42,827)(42,833)(250,833){37}
//: {38}(30,825)(30,803){39}
//: {40}(32,801)(251,801){41}
//: {42}(30,799)(30,764){43}
//: {44}(32,762)(42,762)(42,761)(251,761){45}
//: {46}(30,760)(30,732){47}
//: {48}(32,730)(42,730)(42,729)(252,729){49}
//: {50}(30,728)(30,701){51}
//: {52}(32,699)(42,699)(42,698)(253,698){53}
//: {54}(30,697)(30,668){55}
//: {56}(32,666)(59,666)(59,666)(254,666){57}
//: {58}(30,664)(30,605){59}
//: {60}(32,603)(42,603)(42,601)(253,601){61}
//: {62}(30,601)(30,569){63}
//: {64}(32,567)(42,567)(42,569)(254,569){65}
//: {66}(30,565)(30,541){67}
//: {68}(32,539)(42,539)(42,538)(255,538){69}
//: {70}(30,537)(30,504){71}
//: {72}(32,502)(42,502)(42,506)(256,506){73}
//: {74}(30,500)(30,466){75}
//: {76}(32,464)(42,464)(42,466)(256,466){77}
//: {78}(30,462)(30,436){79}
//: {80}(32,434)(257,434){81}
//: {82}(30,432)(30,402){83}
//: {84}(32,400)(42,400)(42,403)(258,403){85}
//: {86}(30,398)(30,373){87}
//: {88}(32,371)(259,371){89}
//: {90}(30,369)(30,304){91}
//: {92}(32,302)(42,302)(42,301)(256,301){93}
//: {94}(30,300)(30,271){95}
//: {96}(32,269)(257,269){97}
//: {98}(30,267)(30,238){99}
//: {100}(32,236)(42,236)(42,238)(258,238){101}
//: {102}(30,234)(30,208){103}
//: {104}(32,206)(259,206){105}
//: {106}(30,204)(30,168){107}
//: {108}(32,166)(259,166){109}
//: {110}(30,164)(30,137){111}
//: {112}(32,135)(42,135)(42,134)(260,134){113}
//: {114}(30,133)(30,101){115}
//: {116}(32,99)(42,99)(42,101)(256,101){117}
//: {118}(30,97)(30,76){119}
//: {120}(32,74)(42,74)(42,71)(262,71){121}
//: {122}(30,72)(30,19)(97,19)(97,-15){123}
//: {124}(30,1161)(30,1196)(245,1196){125}
wire w97;    //: /sn:0 {0}(245,1191)(73,1191)(73,1159){1}
//: {2}(75,1157)(85,1157)(85,1159)(246,1159){3}
//: {4}(73,1155)(73,1126){5}
//: {6}(75,1124)(85,1124)(85,1128)(247,1128){7}
//: {8}(73,1122)(73,1097){9}
//: {10}(75,1095)(85,1095)(85,1096)(248,1096){11}
//: {12}(73,1093)(73,1057){13}
//: {14}(75,1055)(85,1055)(85,1056)(248,1056){15}
//: {16}(73,1053)(73,1027){17}
//: {18}(75,1025)(85,1025)(85,1024)(249,1024){19}
//: {20}(73,1023)(73,993){21}
//: {22}(75,991)(85,991)(85,993)(250,993){23}
//: {24}(73,989)(73,962){25}
//: {26}(75,960)(85,960)(85,961)(251,961){27}
//: {28}(73,958)(73,894){29}
//: {30}(75,892)(85,892)(85,891)(248,891){31}
//: {32}(73,890)(73,854){33}
//: {34}(75,852)(85,852)(85,859)(249,859){35}
//: {36}(73,850)(73,823){37}
//: {38}(75,821)(85,821)(85,828)(250,828){39}
//: {40}(73,819)(73,798){41}
//: {42}(75,796)(251,796){43}
//: {44}(73,794)(73,754){45}
//: {46}(75,752)(85,752)(85,756)(251,756){47}
//: {48}(73,750)(73,722){49}
//: {50}(75,720)(85,720)(85,724)(252,724){51}
//: {52}(73,718)(73,694){53}
//: {54}(75,692)(85,692)(85,693)(253,693){55}
//: {56}(73,690)(73,664){57}
//: {58}(75,662)(80,662)(80,661)(254,661){59}
//: {60}(73,660)(73,595){61}
//: {62}(75,593)(85,593)(85,596)(253,596){63}
//: {64}(73,591)(73,567){65}
//: {66}(75,565)(85,565)(85,564)(254,564){67}
//: {68}(73,563)(73,539){69}
//: {70}(75,537)(85,537)(85,533)(255,533){71}
//: {72}(73,535)(73,502){73}
//: {74}(75,500)(85,500)(85,501)(256,501){75}
//: {76}(73,498)(73,463){77}
//: {78}(75,461)(256,461){79}
//: {80}(73,459)(73,431){81}
//: {82}(75,429)(257,429){83}
//: {84}(73,427)(73,398){85}
//: {86}(75,396)(85,396)(85,398)(258,398){87}
//: {88}(73,394)(73,364){89}
//: {90}(75,362)(85,362)(85,366)(259,366){91}
//: {92}(73,360)(73,300){93}
//: {94}(75,298)(85,298)(85,296)(256,296){95}
//: {96}(73,296)(73,266){97}
//: {98}(75,264)(257,264){99}
//: {100}(73,262)(73,236){101}
//: {102}(75,234)(85,234)(85,233)(258,233){103}
//: {104}(73,232)(73,198){105}
//: {106}(75,196)(85,196)(85,201)(259,201){107}
//: {108}(73,194)(73,163){109}
//: {110}(75,161)(259,161){111}
//: {112}(73,159)(73,130){113}
//: {114}(75,128)(85,128)(85,129)(260,129){115}
//: {116}(73,126)(73,96){117}
//: {118}(75,94)(85,94)(85,96)(256,96){119}
//: {120}(73,92)(73,70){121}
//: {122}(75,68)(85,68)(85,66)(262,66){123}
//: {124}(73,66)(73,25)(107,25)(107,-15){125}
wire w10;    //: /sn:0 {0}(246,1174)(-51,1174){1}
//: {2}(-53,1172)(-53,1143){3}
//: {4}(-51,1141)(-41,1141)(-41,1143)(247,1143){5}
//: {6}(-53,1139)(-53,1107){7}
//: {8}(-51,1105)(-41,1105)(-41,1111)(248,1111){9}
//: {10}(-53,1103)(-53,1073){11}
//: {12}(-51,1071)(248,1071){13}
//: {14}(-53,1069)(-53,1035){15}
//: {16}(-51,1033)(-41,1033)(-41,1039)(249,1039){17}
//: {18}(-53,1031)(-53,1010){19}
//: {20}(-51,1008)(250,1008){21}
//: {22}(-53,1006)(-53,976){23}
//: {24}(-51,974)(-41,974)(-41,976)(251,976){25}
//: {26}(-53,972)(-53,907){27}
//: {28}(-51,905)(-41,905)(-41,906)(248,906){29}
//: {30}(-53,903)(-53,873){31}
//: {32}(-51,871)(-41,871)(-41,874)(249,874){33}
//: {34}(-53,869)(-53,842){35}
//: {36}(-51,840)(-41,840)(-41,843)(250,843){37}
//: {38}(-53,838)(-53,808){39}
//: {40}(-51,806)(-41,806)(-41,811)(251,811){41}
//: {42}(-53,804)(-53,773){43}
//: {44}(-51,771)(251,771){45}
//: {46}(-53,769)(-53,740){47}
//: {48}(-51,738)(-41,738)(-41,739)(252,739){49}
//: {50}(-53,736)(-53,704){51}
//: {52}(-51,702)(-41,702)(-41,708)(253,708){53}
//: {54}(-53,700)(-53,680){55}
//: {56}(-51,678)(-41,678)(-41,676)(254,676){57}
//: {58}(-53,676)(-53,613){59}
//: {60}(-51,611)(253,611){61}
//: {62}(-53,609)(-53,577){63}
//: {64}(-51,575)(-41,575)(-41,579)(254,579){65}
//: {66}(-53,573)(-53,549){67}
//: {68}(-51,547)(-41,547)(-41,548)(255,548){69}
//: {70}(-53,545)(-53,510){71}
//: {72}(-51,508)(-41,508)(-41,516)(256,516){73}
//: {74}(-53,506)(-53,475){75}
//: {76}(-51,473)(-41,473)(-41,476)(256,476){77}
//: {78}(-53,471)(-53,444){79}
//: {80}(-51,442)(-41,442)(-41,444)(257,444){81}
//: {82}(-53,440)(-53,410){83}
//: {84}(-51,408)(-41,408)(-41,413)(258,413){85}
//: {86}(-53,406)(-53,385){87}
//: {88}(-51,383)(-41,383)(-41,381)(259,381){89}
//: {90}(-53,381)(-53,310){91}
//: {92}(-51,308)(-41,308)(-41,311)(256,311){93}
//: {94}(-53,306)(-53,280){95}
//: {96}(-51,278)(-41,278)(-41,279)(257,279){97}
//: {98}(-53,276)(-53,240){99}
//: {100}(-51,238)(-41,238)(-41,248)(258,248){101}
//: {102}(-53,236)(-53,213){103}
//: {104}(-51,211)(-41,211)(-41,216)(259,216){105}
//: {106}(-53,209)(-53,182){107}
//: {108}(-51,180)(-41,180)(-41,176)(259,176){109}
//: {110}(-53,178)(-53,144){111}
//: {112}(-51,142)(-41,142)(-41,144)(260,144){113}
//: {114}(-53,140)(-53,111){115}
//: {116}(-51,109)(-41,109)(-41,111)(256,111){117}
//: {118}(-53,107)(-53,84){119}
//: {120}(-51,82)(-23,82)(-23,81)(262,81){121}
//: {122}(-53,80)(-53,9)(77,9)(77,-15){123}
//: {124}(-53,1176)(-53,1206)(245,1206){125}
//: enddecls

  //: joint g165 (w4) @(3, 765) /w:[ 44 46 -1 43 ]
  //: joint g154 (w4) @(3, 700) /w:[ 52 54 -1 51 ]
  //: OUT g4 (S3) @(346,166) /sn:0 /w:[ 1 ]
  //: OUT g8 (S7) @(340,302) /sn:0 /w:[ 1 ]
  //: joint g186 (w6) @(117, 955) /w:[ 26 28 -1 25 ]
  //: joint g140 (w10) @(-53, 575) /w:[ 64 66 -1 63 ]
  //: OUT g13 (S12) @(393,488) /sn:0 /w:[ 1 ]
  _GGAND5 #(12) g37 (.I0(w6), .I1(!w97), .I2(w0), .I3(!w4), .I4(!w10), .Z(S5));   //: @(269,238) /sn:0 /w:[ 103 103 101 101 101 0 ]
  _GGAND5 #(12) g55 (.I0(w6), .I1(!w97), .I2(w0), .I3(w4), .I4(w10), .Z(S29));   //: @(258,1133) /sn:0 /w:[ 7 7 5 5 5 0 ]
  _GGAND5 #(12) g58 (.I0(w6), .I1(w97), .I2(!w0), .I3(!w4), .I4(w10), .Z(S19));   //: @(262,761) /sn:0 /w:[ 47 47 45 45 45 0 ]
  //: joint g139 (w4) @(3, 570) /w:[ 64 66 -1 63 ]
  //: joint g112 (w97) @(73, 396) /w:[ 86 88 -1 85 ]
  //: joint g211 (w6) @(117, 1124) /w:[ 6 8 -1 5 ]
  //: joint g76 (w6) @(117, 123) /w:[ 114 116 -1 113 ]
  //: joint g111 (w6) @(117, 393) /w:[ 86 88 -1 85 ]
  //: joint g218 (w0) @(30, 1159) /w:[ 1 2 -1 124 ]
  //: joint g176 (w6) @(117, 852) /w:[ 34 36 -1 33 ]
  //: joint g157 (w97) @(73, 720) /w:[ 50 52 -1 49 ]
  //: joint g163 (w97) @(73, 752) /w:[ 46 48 -1 45 ]
  //: OUT g1 (S0) @(336,74) /sn:0 /w:[ 1 ]
  _GGAND5 #(12) g64 (.I0(!w6), .I1(!w97), .I2(!w0), .I3(!w4), .I4(w10), .Z(S16));   //: @(265,666) /sn:0 /w:[ 59 59 57 57 57 0 ]
  //: joint g166 (w6) @(117, 791) /w:[ 42 44 -1 41 ]
  //: OUT g11 (S10) @(361,446) /sn:0 /w:[ 1 ]
  //: joint g206 (w6) @(117, 1091) /w:[ 10 12 -1 9 ]
  //: joint g130 (w10) @(-53, 508) /w:[ 72 74 -1 71 ]
  //: joint g121 (w97) @(73, 461) /w:[ 78 80 -1 77 ]
  //: OUT g28 (S27) @(369,1067) /sn:0 /w:[ 1 ]
  _GGAND5 #(12) g50 (.I0(w6), .I1(!w97), .I2(w0), .I3(!w4), .I4(w10), .Z(S21));   //: @(261,833) /sn:0 /w:[ 39 39 37 37 37 0 ]
  //: joint g197 (w97) @(73, 1025) /w:[ 18 20 -1 17 ]
  //: joint g132 (w6) @(117, 527) /w:[ 70 72 -1 69 ]
  //: OUT g19 (S18) @(386,737) /sn:0 /w:[ 1 ]
  //: joint g113 (w0) @(30, 400) /w:[ 84 86 -1 83 ]
  //: joint g150 (w10) @(-53, 678) /w:[ 56 58 -1 55 ]
  //: joint g146 (w97) @(73, 662) /w:[ 58 60 -1 57 ]
  //: joint g208 (w0) @(30, 1101) /w:[ 8 10 -1 7 ]
  //: joint g192 (w0) @(30, 998) /w:[ 20 22 -1 19 ]
  //: joint g177 (w0) @(30, 862) /w:[ 32 34 -1 31 ]
  //: OUT g6 (S5) @(339,240) /sn:0 /w:[ 1 ]
  _GGAND5 #(12) g38 (.I0(w6), .I1(w97), .I2(w0), .I3(!w4), .I4(!w10), .Z(S7));   //: @(267,301) /sn:0 /w:[ 95 95 93 93 93 0 ]
  //: joint g115 (w10) @(-53, 408) /w:[ 84 86 -1 83 ]
  //: OUT g7 (S6) @(340,272) /sn:0 /w:[ 1 ]
  _GGAND5 #(12) g53 (.I0(w6), .I1(w97), .I2(w0), .I3(w4), .I4(w10), .Z(S31));   //: @(256,1196) /sn:0 /w:[ 0 0 125 125 125 0 ]
  //: joint g75 (w10) @(-53, 109) /w:[ 116 118 -1 115 ]
  //: joint g169 (w4) @(3, 807) /w:[ 40 42 -1 39 ]
  //: joint g160 (w10) @(-53, 738) /w:[ 48 50 -1 47 ]
  //: joint g135 (w10) @(-53, 547) /w:[ 68 70 -1 67 ]
  //: OUT g20 (S19) @(390,760) /sn:0 /w:[ 1 ]
  //: OUT g31 (S30) @(385,1151) /sn:0 /w:[ 1 ]
  //: joint g149 (w4) @(3, 673) /w:[ 56 58 -1 55 ]
  //: joint g124 (w4) @(3, 470) /w:[ 76 78 -1 75 ]
  //: joint g207 (w97) @(73, 1095) /w:[ 10 12 -1 9 ]
  _GGAND5 #(12) g39 (.I0(!w6), .I1(w97), .I2(w0), .I3(!w4), .I4(!w10), .Z(S6));   //: @(268,269) /sn:0 /w:[ 99 99 97 97 97 0 ]
  //: joint g68 (w0) @(30, 74) /w:[ 120 122 -1 119 ]
  //: joint g200 (w10) @(-53, 1033) /w:[ 16 18 -1 15 ]
  _GGAND5 #(12) g48 (.I0(!w6), .I1(!w97), .I2(!w0), .I3(w4), .I4(!w10), .Z(S8));   //: @(270,371) /sn:0 /w:[ 91 91 89 89 89 0 ]
  //: joint g195 (w10) @(-53, 1008) /w:[ 20 22 -1 19 ]
  //: OUT g17 (S16) @(379,674) /sn:0 /w:[ 1 ]
  //: OUT g25 (S24) @(358,981) /sn:0 /w:[ 1 ]
  //: OUT g29 (S28) @(378,1088) /sn:0 /w:[ 1 ]
  //: joint g205 (w10) @(-53, 1071) /w:[ 12 14 -1 11 ]
  //: joint g179 (w4) @(3, 866) /w:[ 32 34 -1 31 ]
  _GGAND5 #(12) g52 (.I0(!w6), .I1(w97), .I2(w0), .I3(!w4), .I4(w10), .Z(S22));   //: @(260,864) /sn:0 /w:[ 35 35 33 33 33 0 ]
  //: joint g106 (w6) @(117, 359) /w:[ 90 92 -1 89 ]
  //: joint g107 (w0) @(30, 371) /w:[ 88 90 -1 87 ]
  //: joint g174 (w4) @(3, 838) /w:[ 36 38 -1 35 ]
  //: joint g83 (w0) @(30, 166) /w:[ 108 110 -1 107 ]
  //: joint g201 (w6) @(117, 1051) /w:[ 14 16 -1 13 ]
  //: joint g100 (w10) @(-53, 278) /w:[ 96 98 -1 95 ]
  //: OUT g14 (S13) @(382,530) /sn:0 /w:[ 1 ]
  //: joint g202 (w97) @(73, 1055) /w:[ 14 16 -1 13 ]
  //: joint g193 (w97) @(73, 991) /w:[ 22 24 -1 21 ]
  _GGAND5 #(12) g44 (.I0(!w6), .I1(w97), .I2(w0), .I3(w4), .I4(!w10), .Z(S14));   //: @(265,569) /sn:0 /w:[ 67 67 65 65 65 1 ]
  _GGAND5 #(12) g47 (.I0(!w6), .I1(w97), .I2(!w0), .I3(w4), .I4(!w10), .Z(S10));   //: @(268,434) /sn:0 /w:[ 83 83 81 81 81 0 ]
  //: joint g80 (w10) @(-53, 142) /w:[ 112 114 -1 111 ]
  //: joint g94 (w4) @(3, 236) /w:[ 100 102 -1 99 ]
  //: joint g172 (w97) @(73, 821) /w:[ 38 40 -1 37 ]
  //: joint g159 (w4) @(3, 734) /w:[ 48 50 -1 47 ]
  //: OUT g21 (S20) @(356,802) /sn:0 /w:[ 1 ]
  //: joint g84 (w4) @(3, 169) /w:[ 108 110 -1 107 ]
  //: joint g105 (w10) @(-53, 308) /w:[ 92 94 -1 91 ]
  //: joint g155 (w10) @(-53, 702) /w:[ 52 54 -1 51 ]
  //: joint g141 (w6) @(117, 586) /w:[ 62 64 -1 61 ]
  //: OUT g23 (S22) @(363,865) /sn:0 /w:[ 1 ]
  _GGAND5 #(12) g41 (.I0(w6), .I1(!w97), .I2(!w0), .I3(w4), .I4(!w10), .Z(S9));   //: @(269,403) /sn:0 /w:[ 87 87 85 85 85 0 ]
  //: joint g151 (w6) @(117, 687) /w:[ 54 56 -1 53 ]
  _GGAND5 #(12) g40 (.I0(!w6), .I1(!w97), .I2(w0), .I3(!w4), .I4(!w10), .Z(S4));   //: @(270,206) /sn:0 /w:[ 107 107 105 105 105 1 ]
  _GGAND5 #(12) g54 (.I0(!w6), .I1(!w97), .I2(!w0), .I3(w4), .I4(w10), .Z(S24));   //: @(262,966) /sn:0 /w:[ 27 27 25 25 25 0 ]
  //: joint g93 (w0) @(30, 236) /w:[ 100 102 -1 99 ]
  //: joint g116 (w6) @(117, 426) /w:[ 82 84 -1 81 ]
  //: joint g123 (w0) @(30, 464) /w:[ 76 78 -1 75 ]
  //: joint g167 (w97) @(73, 796) /w:[ 42 44 -1 41 ]
  //: IN g0 (C) @(94,-108) /sn:0 /R:3 /w:[ 1 ]
  //: OUT g26 (S25) @(359,1006) /sn:0 /w:[ 1 ]
  _GGAND5 #(12) g46 (.I0(!w6), .I1(!w97), .I2(w0), .I3(w4), .I4(!w10), .Z(S12));   //: @(267,506) /sn:0 /w:[ 75 75 73 73 73 0 ]
  //: joint g90 (w10) @(-53, 211) /w:[ 104 106 -1 103 ]
  //: joint g82 (w97) @(73, 161) /w:[ 110 112 -1 109 ]
  //: joint g136 (w6) @(117, 556) /w:[ 66 68 -1 65 ]
  //: joint g128 (w4) @(3, 508) /w:[ 72 74 -1 71 ]
  //: joint g190 (w10) @(-53, 974) /w:[ 24 26 -1 23 ]
  //: joint g173 (w0) @(30, 827) /w:[ 36 38 -1 35 ]
  _GGAND5 #(10) g33 (.I0(!w6), .I1(!w97), .I2(!w0), .I3(!w4), .I4(!w10), .Z(S0));   //: @(273,71) /sn:0 /w:[ 123 123 121 121 121 0 ]
  //: joint g91 (w97) @(73, 234) /w:[ 102 104 -1 101 ]
  _GGAND5 #(12) g49 (.I0(w6), .I1(!w97), .I2(!w0), .I3(!w4), .I4(w10), .Z(S17));   //: @(264,698) /sn:0 /w:[ 55 55 53 53 53 0 ]
  //: joint g198 (w0) @(30, 1023) /w:[ 16 18 -1 15 ]
  //: joint g137 (w97) @(73, 565) /w:[ 66 68 -1 65 ]
  _GGAND5 #(12) g61 (.I0(!w6), .I1(w97), .I2(!w0), .I3(!w4), .I4(w10), .Z(S18));   //: @(263,729) /sn:0 /w:[ 51 51 49 49 49 0 ]
  //: joint g220 (w4) @(3, 1168) /w:[ 1 2 -1 124 ]
  //: joint g158 (w0) @(30, 730) /w:[ 48 50 -1 47 ]
  //: OUT g3 (S2) @(340,140) /sn:0 /w:[ 0 ]
  _GGAND5 #(12) g34 (.I0(w6), .I1(!w97), .I2(!w0), .I3(!w4), .I4(!w10), .Z(S1));   //: @(267,101) /sn:0 /w:[ 119 119 117 117 117 0 ]
  _GGAND5 #(12) g51 (.I0(w6), .I1(w97), .I2(w0), .I3(!w4), .I4(w10), .Z(S23));   //: @(259,896) /sn:0 /w:[ 31 31 29 29 29 0 ]
  //: joint g86 (w6) @(117, 193) /w:[ 106 108 -1 105 ]
  //: joint g217 (w97) @(73, 1157) /w:[ 2 4 -1 1 ]
  //: joint g89 (w4) @(3, 208) /w:[ 104 106 -1 103 ]
  //: OUT g2 (S1) @(342,104) /sn:0 /w:[ 1 ]
  assign {w10, w4, w0, w97, w6} = C; //: CONCAT g65  @(97,-20) /sn:0 /R:1 /w:[ 123 123 123 125 125 0 ] /dr:0 /tp:0 /drp:0
  //: joint g77 (w97) @(73, 128) /w:[ 114 116 -1 113 ]
  //: joint g110 (w10) @(-53, 383) /w:[ 88 90 -1 87 ]
  //: joint g213 (w0) @(30, 1130) /w:[ 4 6 -1 3 ]
  //: joint g156 (w6) @(117, 717) /w:[ 50 52 -1 49 ]
  //: joint g148 (w0) @(30, 666) /w:[ 56 58 -1 55 ]
  //: joint g147 (w6) @(117, 647) /w:[ 58 60 -1 57 ]
  _GGAND5 #(12) g59 (.I0(w6), .I1(!w97), .I2(!w0), .I3(w4), .I4(w10), .Z(S25));   //: @(261,998) /sn:0 /w:[ 23 23 21 21 21 0 ]
  //: joint g203 (w0) @(30, 1060) /w:[ 12 14 -1 11 ]
  //: joint g153 (w97) @(73, 692) /w:[ 54 56 -1 53 ]
  //: joint g72 (w97) @(73, 94) /w:[ 118 120 -1 117 ]
  //: joint g196 (w6) @(117, 1020) /w:[ 18 20 -1 17 ]
  //: joint g182 (w97) @(73, 892) /w:[ 30 32 -1 29 ]
  //: joint g161 (w6) @(117, 752) /w:[ 46 48 -1 45 ]
  //: joint g98 (w0) @(30, 269) /w:[ 96 98 -1 95 ]
  //: joint g99 (w4) @(3, 274) /w:[ 96 98 -1 95 ]
  //: OUT g16 (S15) @(404,574) /sn:0 /w:[ 0 ]
  //: joint g96 (w6) @(117, 259) /w:[ 98 100 -1 97 ]
  //: joint g189 (w4) @(3, 969) /w:[ 24 26 -1 23 ]
  //: joint g183 (w0) @(30, 894) /w:[ 28 30 -1 27 ]
  //: joint g152 (w0) @(30, 699) /w:[ 52 54 -1 51 ]
  //: joint g103 (w0) @(30, 302) /w:[ 92 94 -1 91 ]
  //: joint g122 (w6) @(117, 454) /w:[ 78 80 -1 77 ]
  //: joint g212 (w97) @(73, 1124) /w:[ 6 8 -1 5 ]
  //: OUT g10 (S9) @(355,408) /sn:0 /w:[ 1 ]
  //: joint g78 (w0) @(30, 135) /w:[ 112 114 -1 111 ]
  //: joint g87 (w97) @(73, 196) /w:[ 106 108 -1 105 ]
  //: joint g199 (w4) @(3, 1028) /w:[ 16 18 -1 15 ]
  //: joint g171 (w6) @(117, 823) /w:[ 38 40 -1 37 ]
  //: joint g129 (w0) @(30, 502) /w:[ 72 74 -1 71 ]
  //: OUT g27 (S26) @(365,1044) /sn:0 /w:[ 1 ]
  //: OUT g32 (S31) @(350,1211) /sn:0 /w:[ 1 ]
  //: joint g187 (w0) @(30, 964) /w:[ 24 26 -1 23 ]
  //: joint g102 (w97) @(73, 298) /w:[ 94 96 -1 93 ]
  //: joint g143 (w0) @(30, 603) /w:[ 60 62 -1 59 ]
  //: joint g69 (w4) @(3, 76) /w:[ 120 122 -1 119 ]
  //: OUT g9 (S8) @(354,383) /sn:0 /w:[ 1 ]
  _GGAND5 #(12) g57 (.I0(!w6), .I1(w97), .I2(!w0), .I3(w4), .I4(w10), .Z(S26));   //: @(260,1029) /sn:0 /w:[ 19 19 17 17 17 0 ]
  //: joint g119 (w4) @(3, 440) /w:[ 80 82 -1 79 ]
  //: joint g142 (w97) @(73, 593) /w:[ 62 64 -1 61 ]
  //: OUT g15 (S14) @(400,551) /sn:0 /w:[ 0 ]
  //: joint g71 (w6) @(117, 92) /w:[ 118 120 -1 117 ]
  //: joint g162 (w0) @(30, 762) /w:[ 44 46 -1 43 ]
  //: joint g131 (w97) @(73, 537) /w:[ 70 72 -1 69 ]
  //: joint g67 (w97) @(73, 68) /w:[ 122 124 -1 121 ]
  //: joint g127 (w97) @(73, 500) /w:[ 74 76 -1 73 ]
  _GGAND5 #(12) g43 (.I0(w6), .I1(w97), .I2(w0), .I3(w4), .I4(!w10), .Z(S15));   //: @(264,601) /sn:0 /w:[ 63 63 61 61 61 1 ]
  //: joint g145 (w10) @(-53, 611) /w:[ 60 62 -1 59 ]
  _GGAND5 #(12) g62 (.I0(w6), .I1(w97), .I2(!w0), .I3(w4), .I4(w10), .Z(S27));   //: @(259,1061) /sn:0 /w:[ 15 15 13 13 13 0 ]
  //: joint g73 (w0) @(30, 99) /w:[ 116 118 -1 115 ]
  //: joint g88 (w0) @(30, 206) /w:[ 104 106 -1 103 ]
  //: joint g104 (w4) @(3, 306) /w:[ 92 94 -1 91 ]
  //: joint g188 (w97) @(73, 960) /w:[ 26 28 -1 25 ]
  //: joint g180 (w10) @(-53, 871) /w:[ 32 34 -1 31 ]
  //: joint g138 (w0) @(30, 567) /w:[ 64 66 -1 63 ]
  _GGAND5 #(12) g42 (.I0(w6), .I1(!w97), .I2(w0), .I3(w4), .I4(!w10), .Z(S13));   //: @(266,538) /sn:0 /w:[ 71 71 69 69 69 0 ]
  _GGAND5 #(12) g63 (.I0(!w6), .I1(!w97), .I2(w0), .I3(w4), .I4(w10), .Z(S28));   //: @(259,1101) /sn:0 /w:[ 11 11 9 9 9 0 ]
  //: joint g175 (w10) @(-53, 840) /w:[ 36 38 -1 35 ]
  //: joint g74 (w4) @(3, 104) /w:[ 116 118 -1 115 ]
  //: joint g109 (w4) @(3, 375) /w:[ 88 90 -1 87 ]
  //: joint g181 (w6) @(117, 885) /w:[ 30 32 -1 29 ]
  //: joint g168 (w0) @(30, 801) /w:[ 40 42 -1 39 ]
  //: joint g133 (w0) @(30, 539) /w:[ 68 70 -1 67 ]
  //: OUT g5 (S4) @(336,207) /sn:0 /w:[ 0 ]
  _GGAND5 #(12) g56 (.I0(!w6), .I1(w97), .I2(w0), .I3(w4), .I4(w10), .Z(S30));   //: @(257,1164) /sn:0 /w:[ 3 3 0 0 0 0 ]
  //: joint g215 (w10) @(-53, 1141) /w:[ 4 6 -1 3 ]
  //: joint g194 (w4) @(3, 1002) /w:[ 20 22 -1 19 ]
  //: joint g79 (w4) @(3, 138) /w:[ 112 114 -1 111 ]
  //: joint g95 (w10) @(-53, 238) /w:[ 100 102 -1 99 ]
  //: joint g117 (w97) @(73, 429) /w:[ 82 84 -1 81 ]
  //: joint g216 (w6) @(117, 1151) /w:[ 2 4 -1 1 ]
  //: OUT g24 (S23) @(367,888) /sn:0 /w:[ 1 ]
  _GGAND5 #(12) g36 (.I0(w6), .I1(w97), .I2(!w0), .I3(!w4), .I4(!w10), .Z(S3));   //: @(270,166) /sn:0 /w:[ 111 111 109 109 109 0 ]
  //: joint g85 (w10) @(-53, 180) /w:[ 108 110 -1 107 ]
  //: joint g92 (w6) @(117, 228) /w:[ 102 104 -1 101 ]
  //: joint g178 (w97) @(73, 852) /w:[ 34 36 -1 33 ]
  //: joint g144 (w4) @(3, 606) /w:[ 60 62 -1 59 ]
  //: joint g125 (w10) @(-53, 473) /w:[ 76 78 -1 75 ]
  //: joint g214 (w4) @(3, 1135) /w:[ 4 6 -1 3 ]
  //: joint g210 (w10) @(-53, 1105) /w:[ 8 10 -1 7 ]
  _GGAND5 #(12) g60 (.I0(!w6), .I1(!w97), .I2(w0), .I3(!w4), .I4(w10), .Z(S20));   //: @(262,801) /sn:0 /w:[ 43 43 41 41 41 0 ]
  //: joint g81 (w6) @(117, 156) /w:[ 110 112 -1 109 ]
  //: joint g101 (w6) @(117, 292) /w:[ 94 96 -1 93 ]
  //: joint g204 (w4) @(3, 1064) /w:[ 12 14 -1 11 ]
  //: joint g185 (w10) @(-53, 905) /w:[ 28 30 -1 27 ]
  //: joint g170 (w10) @(-53, 806) /w:[ 40 42 -1 39 ]
  //: OUT g22 (S21) @(357,827) /sn:0 /w:[ 1 ]
  _GGAND5 #(12) g35 (.I0(!w6), .I1(w97), .I2(!w0), .I3(!w4), .I4(!w10), .Z(S2));   //: @(271,134) /sn:0 /w:[ 115 115 113 113 113 1 ]
  _GGAND5 #(12) g45 (.I0(w6), .I1(w97), .I2(!w0), .I3(w4), .I4(!w10), .Z(S11));   //: @(267,466) /sn:0 /w:[ 79 79 77 77 77 0 ]
  //: joint g70 (w10) @(-53, 82) /w:[ 120 122 -1 119 ]
  //: joint g126 (w6) @(117, 496) /w:[ 74 76 -1 73 ]
  //: joint g209 (w4) @(3, 1106) /w:[ 8 10 -1 7 ]
  //: joint g184 (w4) @(3, 900) /w:[ 28 30 -1 27 ]
  //: joint g66 (w6) @(117, 62) /w:[ 122 124 -1 121 ]
  //: joint g97 (w97) @(73, 264) /w:[ 98 100 -1 97 ]
  //: joint g114 (w4) @(3, 406) /w:[ 84 86 -1 83 ]
  //: joint g120 (w10) @(-53, 442) /w:[ 80 82 -1 79 ]
  //: OUT g12 (S11) @(365,469) /sn:0 /w:[ 1 ]
  //: OUT g18 (S17) @(380,699) /sn:0 /w:[ 1 ]
  //: joint g219 (w10) @(-53, 1174) /w:[ 1 2 -1 124 ]
  //: joint g191 (w6) @(117, 988) /w:[ 22 24 -1 21 ]
  //: joint g164 (w10) @(-53, 771) /w:[ 44 46 -1 43 ]
  //: OUT g30 (S29) @(379,1113) /sn:0 /w:[ 1 ]
  //: joint g108 (w97) @(73, 362) /w:[ 90 92 -1 89 ]
  //: joint g134 (w4) @(3, 542) /w:[ 68 70 -1 67 ]
  //: joint g118 (w0) @(30, 434) /w:[ 80 82 -1 79 ]

endmodule
//: /netlistEnd

//: /netlistBegin Banco32Reg
module Banco32Reg(Leer1, Reloj, RegLeer1, RegEsc, Leer2, W, Esc, RegLeer2);
//: interface  /sz:(128, 112) /bd:[ Ti0>W(61/128) Li0>RegLeer2[4:0](38/112) Li1>RegLeer1[4:0](17/112) Li2>RegEsc[4:0](63/112) Li3>Esc[31:0](85/112) Bi0>Reloj(64/128) Ro0<Leer2[31:0](72/112) Ro1<Leer1[31:0](37/112) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [4:0] RegEsc;    //: /sn:0 {0}(#:-279,700)(-150,700)(-150,699)(#:-146,699){1}
output [31:0] Leer1;    //: /sn:0 {0}(#:1266,627)(1196,627)(1196,713)(1011,713)(1011,696)(993,696){1}
input [31:0] Esc;    //: /sn:0 {0}(#:457,1348)(377,1348)(377,1353)(367,1353){1}
//: {2}(365,1351)(365,1311){3}
//: {4}(367,1309)(377,1309)(377,1307)(#:457,1307){5}
//: {6}(365,1307)(365,1269){7}
//: {8}(367,1267)(377,1267)(377,1266)(#:457,1266){9}
//: {10}(365,1265)(365,1229){11}
//: {12}(367,1227)(377,1227)(377,1225)(#:457,1225){13}
//: {14}(365,1225)(365,1188){15}
//: {16}(367,1186)(377,1186)(377,1184)(#:457,1184){17}
//: {18}(365,1184)(365,1145){19}
//: {20}(367,1143)(#:457,1143){21}
//: {22}(365,1141)(365,1104){23}
//: {24}(367,1102)(#:457,1102){25}
//: {26}(365,1100)(365,1062){27}
//: {28}(367,1060)(377,1060)(377,1061)(#:457,1061){29}
//: {30}(365,1058)(365,1007){31}
//: {32}(367,1005)(#:458,1005){33}
//: {34}(365,1003)(365,969){35}
//: {36}(367,967)(377,967)(377,964)(#:458,964){37}
//: {38}(365,965)(365,924){39}
//: {40}(367,922)(377,922)(377,923)(#:458,923){41}
//: {42}(365,920)(365,884){43}
//: {44}(367,882)(#:458,882){45}
//: {46}(365,880)(365,844){47}
//: {48}(367,842)(377,842)(377,841)(#:458,841){49}
//: {50}(365,840)(365,802){51}
//: {52}(367,800)(#:458,800){53}
//: {54}(365,798)(365,765){55}
//: {56}(367,763)(377,763)(377,759)(#:458,759){57}
//: {58}(365,761)(365,720){59}
//: {60}(367,718)(#:458,718){61}
//: {62}(365,716)(365,663){63}
//: {64}(367,661)(#:457,661){65}
//: {66}(365,659)(365,626){67}
//: {68}(367,624)(377,624)(377,620)(#:457,620){69}
//: {70}(365,622)(365,581){71}
//: {72}(367,579)(#:457,579){73}
//: {74}(365,577)(365,538){75}
//: {76}(367,536)(377,536)(377,538)(#:457,538){77}
//: {78}(365,534)(365,497){79}
//: {80}(367,495)(377,495)(377,497)(#:457,497){81}
//: {82}(365,493)(365,457){83}
//: {84}(367,455)(377,455)(377,456)(#:457,456){85}
//: {86}(365,453)(365,417){87}
//: {88}(367,415)(#:457,415){89}
//: {90}(365,413)(365,373){91}
//: {92}(367,371)(377,371)(377,374)(#:457,374){93}
//: {94}(365,369)(365,313){95}
//: {96}(367,311)(377,311)(377,313)(#:455,313){97}
//: {98}(365,309)(365,274){99}
//: {100}(367,272)(#:455,272){101}
//: {102}(365,270)(365,229){103}
//: {104}(367,227)(377,227)(377,231)(#:455,231){105}
//: {106}(365,225)(365,191){107}
//: {108}(367,189)(377,189)(377,190)(#:455,190){109}
//: {110}(365,187)(365,150){111}
//: {112}(367,148)(377,148)(377,149)(#:455,149){113}
//: {114}(365,146)(365,109){115}
//: {116}(367,107)(377,107)(377,108)(#:455,108){117}
//: {118}(365,105)(365,69){119}
//: {120}(367,67)(#:455,67){121}
//: {122}(365,65)(365,26)(#:455,26){123}
//: {124}(365,1355)(365,1422)(#:326,1422){125}
input [4:0] RegLeer2;    //: /sn:0 {0}(#:1147,282)(1157,282)(1157,297)(1122,297)(1122,328){1}
input Reloj;    //: /sn:0 {0}(457,1358)(425,1358)(425,1357)(415,1357){1}
//: {2}(413,1355)(413,1318){3}
//: {4}(415,1316)(425,1316)(425,1317)(457,1317){5}
//: {6}(413,1314)(413,1279){7}
//: {8}(415,1277)(425,1277)(425,1276)(457,1276){9}
//: {10}(413,1275)(413,1237){11}
//: {12}(415,1235)(457,1235){13}
//: {14}(413,1233)(413,1193){15}
//: {16}(415,1191)(425,1191)(425,1194)(457,1194){17}
//: {18}(413,1189)(413,1155){19}
//: {20}(415,1153)(457,1153){21}
//: {22}(413,1151)(413,1114){23}
//: {24}(415,1112)(457,1112){25}
//: {26}(413,1110)(413,1075){27}
//: {28}(415,1073)(425,1073)(425,1071)(457,1071){29}
//: {30}(413,1071)(413,1014){31}
//: {32}(415,1012)(425,1012)(425,1015)(458,1015){33}
//: {34}(413,1010)(413,977){35}
//: {36}(415,975)(425,975)(425,974)(458,974){37}
//: {38}(413,973)(413,936){39}
//: {40}(415,934)(425,934)(425,933)(458,933){41}
//: {42}(413,932)(413,894){43}
//: {44}(415,892)(458,892){45}
//: {46}(413,890)(413,852){47}
//: {48}(415,850)(425,850)(425,851)(458,851){49}
//: {50}(413,848)(413,813){51}
//: {52}(415,811)(425,811)(425,810)(458,810){53}
//: {54}(413,809)(413,772){55}
//: {56}(415,770)(425,770)(425,769)(458,769){57}
//: {58}(413,768)(413,734){59}
//: {60}(415,732)(425,732)(425,728)(458,728){61}
//: {62}(413,730)(413,672){63}
//: {64}(415,670)(425,670)(425,671)(457,671){65}
//: {66}(413,668)(413,630){67}
//: {68}(415,628)(425,628)(425,630)(457,630){69}
//: {70}(413,626)(413,591){71}
//: {72}(415,589)(457,589){73}
//: {74}(413,587)(413,550){75}
//: {76}(415,548)(457,548){77}
//: {78}(413,546)(413,509){79}
//: {80}(415,507)(457,507){81}
//: {82}(413,505)(413,466){83}
//: {84}(415,464)(425,464)(425,466)(457,466){85}
//: {86}(413,462)(413,425){87}
//: {88}(415,423)(425,423)(425,425)(457,425){89}
//: {90}(413,421)(413,386){91}
//: {92}(415,384)(457,384){93}
//: {94}(413,382)(413,325){95}
//: {96}(415,323)(455,323){97}
//: {98}(413,321)(413,284){99}
//: {100}(415,282)(455,282){101}
//: {102}(413,280)(413,246){103}
//: {104}(415,244)(425,244)(425,241)(455,241){105}
//: {106}(413,242)(413,204){107}
//: {108}(415,202)(425,202)(425,200)(455,200){109}
//: {110}(413,200)(413,163){111}
//: {112}(415,161)(425,161)(425,159)(455,159){113}
//: {114}(413,159)(413,118){115}
//: {116}(415,116)(425,116)(425,118)(455,118){117}
//: {118}(413,114)(413,77){119}
//: {120}(415,75)(425,75)(425,77)(455,77){121}
//: {122}(413,73)(413,36)(455,36){123}
//: {124}(413,1359)(413,1477)(337,1477){125}
input W;    //: /sn:0 {0}(-141,203)(-56,203)(-56,285){1}
//: {2}(-54,287)(-15,287){3}
//: {4}(-56,289)(-56,311){5}
//: {6}(-54,313)(-44,313)(-44,315)(-15,315){7}
//: {8}(-56,315)(-56,343){9}
//: {10}(-54,345)(-44,345)(-44,344)(-15,344){11}
//: {12}(-56,347)(-56,375){13}
//: {14}(-54,377)(-44,377)(-44,373)(-15,373){15}
//: {16}(-56,379)(-56,408){17}
//: {18}(-54,410)(-44,410)(-44,403)(-15,403){19}
//: {20}(-56,412)(-56,437){21}
//: {22}(-54,439)(-44,439)(-44,431)(-15,431){23}
//: {24}(-56,441)(-56,462){25}
//: {26}(-54,464)(-44,464)(-44,460)(-15,460){27}
//: {28}(-56,466)(-56,489){29}
//: {30}(-54,491)(-44,491)(-44,488)(-15,488){31}
//: {32}(-56,493)(-56,519){33}
//: {34}(-54,521)(-44,521)(-44,520)(-13,520){35}
//: {36}(-56,523)(-56,551){37}
//: {38}(-54,553)(-44,553)(-44,548)(-13,548){39}
//: {40}(-56,555)(-56,579){41}
//: {42}(-54,581)(-44,581)(-44,577)(-13,577){43}
//: {44}(-56,583)(-56,610){45}
//: {46}(-54,612)(-44,612)(-44,606)(-13,606){47}
//: {48}(-56,614)(-56,638){49}
//: {50}(-54,640)(-44,640)(-44,636)(-13,636){51}
//: {52}(-56,642)(-56,667){53}
//: {54}(-54,669)(-44,669)(-44,664)(-13,664){55}
//: {56}(-56,671)(-56,696){57}
//: {58}(-54,698)(-44,698)(-44,693)(-13,693){59}
//: {60}(-56,700)(-56,723){61}
//: {62}(-54,725)(-44,725)(-44,721)(-13,721){63}
//: {64}(-56,727)(-56,750){65}
//: {66}(-54,752)(-15,752){67}
//: {68}(-56,754)(-56,784){69}
//: {70}(-54,786)(-44,786)(-44,780)(-15,780){71}
//: {72}(-56,788)(-56,817){73}
//: {74}(-54,819)(-44,819)(-44,809)(-15,809){75}
//: {76}(-56,821)(-56,841){77}
//: {78}(-54,843)(-44,843)(-44,838)(-15,838){79}
//: {80}(-56,845)(-56,872){81}
//: {82}(-54,874)(-44,874)(-44,868)(-15,868){83}
//: {84}(-56,876)(-56,901){85}
//: {86}(-54,903)(-44,903)(-44,896)(-15,896){87}
//: {88}(-56,905)(-56,928){89}
//: {90}(-54,930)(-44,930)(-44,925)(-15,925){91}
//: {92}(-56,932)(-56,957){93}
//: {94}(-54,959)(-44,959)(-44,953)(-15,953){95}
//: {96}(-56,961)(-56,990){97}
//: {98}(-54,992)(-44,992)(-44,986)(-12,986){99}
//: {100}(-56,994)(-56,1020){101}
//: {102}(-54,1022)(-44,1022)(-44,1014)(-12,1014){103}
//: {104}(-56,1024)(-56,1045){105}
//: {106}(-54,1047)(-44,1047)(-44,1043)(-12,1043){107}
//: {108}(-56,1049)(-56,1078){109}
//: {110}(-54,1080)(-44,1080)(-44,1072)(-12,1072){111}
//: {112}(-56,1082)(-56,1103){113}
//: {114}(-54,1105)(-44,1105)(-44,1102)(-12,1102){115}
//: {116}(-56,1107)(-56,1132){117}
//: {118}(-54,1134)(-44,1134)(-44,1130)(-12,1130){119}
//: {120}(-56,1136)(-56,1160){121}
//: {122}(-54,1162)(-44,1162)(-44,1159)(-12,1159){123}
//: {124}(-56,1164)(-56,1187)(-12,1187){125}
input [4:0] RegLeer1;    //: /sn:0 {0}(#:1006,284)(1016,284)(1016,299)(971,299)(971,337){1}
output [31:0] Leer2;    //: /sn:0 {0}(#:1144,687)(1266,687){1}
wire w160;    //: /sn:0 {0}(-104,281)(-30,281)(-30,282)(-15,282){1}
wire [31:0] w7;    //: /sn:0 {0}(#:586,76)(927,76)(927,387)(937,387){1}
//: {2}(941,387)(951,387){3}
//: {4}(#:939,385)(939,378)(1102,378){5}
wire [31:0] w99;    //: /sn:0 {0}(#:588,1234)(750,1234)(750,1050)(935,1050){1}
//: {2}(939,1050)(951,1050){3}
//: {4}(#:937,1048)(937,1041)(1102,1041){5}
wire w122;    //: /sn:0 {0}(457,1327)(30,1327)(30,1157)(9,1157){1}
wire w134;    //: /sn:0 {0}(-104,1035)(-27,1035)(-27,1038)(-12,1038){1}
wire [31:0] w203;    //: /sn:0 {0}(#:588,1070)(697,1070)(697,951)(935,951){1}
//: {2}(939,951)(#:951,951){3}
//: {4}(#:937,949)(937,942)(1102,942){5}
wire w46;    //: /sn:0 {0}(8,546)(114,546)(114,435)(457,435){1}
wire w135;    //: /sn:0 {0}(-104,1006)(-27,1006)(-27,1009)(-12,1009){1}
wire w153;    //: /sn:0 {0}(-104,484)(-30,484)(-30,483)(-15,483){1}
wire w141;    //: /sn:0 {0}(-104,832)(-30,832)(-30,833)(-15,833){1}
wire [31:0] w19;    //: /sn:0 {0}(#:586,281)(887,281)(887,509)(934,509){1}
//: {2}(938,509)(951,509){3}
//: {4}(#:936,507)(936,500)(1102,500){5}
wire w4;    //: /sn:0 {0}(6,313)(51,313)(51,87)(455,87){1}
wire [31:0] w15;    //: /sn:0 {0}(#:586,117)(920,117)(920,411)(938,411){1}
//: {2}(942,411)(951,411){3}
//: {4}(#:940,409)(940,402)(1102,402){5}
wire w38;    //: /sn:0 {0}(8,575)(120,575)(120,476)(457,476){1}
wire w106;    //: /sn:0 {0}(457,1204)(50,1204)(50,1070)(9,1070){1}
wire [31:0] w51;    //: /sn:0 {0}(#:588,670)(818,670)(818,730)(932,730){1}
//: {2}(936,730)(951,730){3}
//: {4}(#:934,728)(934,721)(1102,721){5}
wire w152;    //: /sn:0 {0}(-104,513)(-28,513)(-28,515)(-13,515){1}
wire w129;    //: /sn:0 {0}(-104,1180)(-27,1180)(-27,1182)(-12,1182){1}
wire w0;    //: /sn:0 {0}(6,285)(44,285)(44,46)(455,46){1}
wire w151;    //: /sn:0 {0}(-104,542)(-28,542)(-28,543)(-13,543){1}
wire w114;    //: /sn:0 {0}(457,1368)(24,1368)(24,1185)(9,1185){1}
wire w66;    //: /sn:0 {0}(458,902)(101,902)(101,866)(6,866){1}
wire [31:0] w111;    //: /sn:0 {0}(#:588,1111)(710,1111)(710,976)(933,976){1}
//: {2}(937,976)(951,976){3}
//: {4}(#:935,974)(935,967)(1102,967){5}
wire w34;    //: /sn:0 {0}(8,634)(134,634)(134,558)(457,558){1}
wire w133;    //: /sn:0 {0}(-104,1064)(-27,1064)(-27,1067)(-12,1067){1}
wire [31:0] w63;    //: /sn:0 {0}(#:588,383)(872,383)(872,559)(935,559){1}
//: {2}(939,559)(951,559){3}
//: {4}(#:937,557)(937,550)(1102,550){5}
wire w159;    //: /sn:0 {0}(-104,310)(-15,310){1}
wire w102;    //: /sn:0 {0}(457,1163)(57,1163)(57,1041)(9,1041){1}
wire [31:0] w87;    //: /sn:0 {0}(#:589,932)(645,932)(645,878)(934,878){1}
//: {2}(938,878)(951,878){3}
//: {4}(#:936,876)(936,869)(1102,869){5}
wire [31:0] w43;    //: /sn:0 {0}(#:588,506)(848,506)(848,632)(935,632){1}
//: {2}(939,632)(951,632){3}
//: {4}(#:937,630)(937,623)(1102,623){5}
wire w157;    //: /sn:0 {0}(-104,368)(-15,368){1}
wire [31:0] w75;    //: /sn:0 {0}(#:951,829)(939,829){1}
//: {2}(#:937,827)(937,820)(1102,820){3}
//: {4}(935,829)(602,829)(#:602,850)(#:589,850){5}
wire [31:0] w119;    //: /sn:0 {0}(#:588,1275)(779,1275)(779,1074)(934,1074){1}
//: {2}(938,1074)(951,1074){3}
//: {4}(#:936,1072)(936,1065)(1102,1065){5}
wire [31:0] w67;    //: /sn:0 {0}(#:951,853)(941,853){1}
//: {2}(#:939,851)(939,844)(1102,844){3}
//: {4}(937,853)(622,853)(#:622,891)(#:589,891){5}
wire w54;    //: /sn:0 {0}(8,662)(141,662)(141,599)(457,599){1}
wire w90;    //: /sn:0 {0}(458,984)(88,984)(88,923)(6,923){1}
wire w58;    //: /sn:0 {0}(8,691)(147,691)(147,640)(457,640){1}
wire [31:0] w31;    //: /sn:0 {0}(#:586,199)(904,199)(904,460)(937,460){1}
//: {2}(941,460)(951,460){3}
//: {4}(#:939,458)(939,451)(1102,451){5}
wire w130;    //: /sn:0 {0}(-104,1151)(-27,1151)(-27,1154)(-12,1154){1}
wire w156;    //: /sn:0 {0}(-104,397)(-30,397)(-30,398)(-15,398){1}
wire [31:0] w23;    //: /sn:0 {0}(#:586,322)(880,322)(880,534)(933,534){1}
//: {2}(937,534)(951,534){3}
//: {4}(#:935,532)(935,525)(1102,525){5}
wire w132;    //: /sn:0 {0}(-104,1093)(-27,1093)(-27,1097)(-12,1097){1}
wire w140;    //: /sn:0 {0}(-104,861)(-30,861)(-30,863)(-15,863){1}
wire w126;    //: /sn:0 {0}(457,1081)(73,1081)(73,984)(9,984){1}
wire w82;    //: /sn:0 {0}(458,1025)(80,1025)(80,951)(6,951){1}
wire w154;    //: /sn:0 {0}(-104,455)(-15,455){1}
wire w74;    //: /sn:0 {0}(6,836)(108,836)(108,861)(458,861){1}
wire w158;    //: /sn:0 {0}(-104,339)(-15,339){1}
wire w98;    //: /sn:0 {0}(9,1100)(42,1100)(42,1245)(457,1245){1}
wire [31:0] w103;    //: /sn:0 {0}(#:588,1152)(721,1152)(721,1001)(932,1001){1}
//: {2}(936,1001)(951,1001){3}
//: {4}(#:934,999)(934,992)(1102,992){5}
wire w8;    //: /sn:0 {0}(6,371)(66,371)(66,169)(455,169){1}
wire [31:0] w91;    //: /sn:0 {0}(#:589,973)(668,973)(668,902)(935,902){1}
//: {2}(939,902)(951,902){3}
//: {4}(#:937,900)(937,893)(1102,893){5}
wire [31:0] w35;    //: /sn:0 {0}(#:588,547)(840,547)(840,657)(936,657){1}
//: {2}(940,657)(951,657){3}
//: {4}(#:938,655)(938,648)(1102,648){5}
wire w118;    //: /sn:0 {0}(457,1286)(35,1286)(35,1128)(9,1128){1}
wire w18;    //: /sn:0 {0}(6,458)(91,458)(91,292)(455,292){1}
wire [31:0] w71;    //: /sn:0 {0}(#:589,809)(660,809)(660,804)(934,804){1}
//: {2}(938,804)(951,804){3}
//: {4}(#:936,802)(936,795)(1102,795){5}
wire w30;    //: /sn:0 {0}(6,401)(75,401)(75,210)(455,210){1}
wire w146;    //: /sn:0 {0}(-104,687)(-28,687)(-28,688)(-13,688){1}
wire w149;    //: /sn:0 {0}(-104,600)(-28,600)(-28,601)(-13,601){1}
wire w22;    //: /sn:0 {0}(6,486)(99,486)(99,333)(455,333){1}
wire w144;    //: /sn:0 {0}(-104,745)(-30,745)(-30,747)(-15,747){1}
wire [31:0] w123;    //: /sn:0 {0}(#:588,1316)(816,1316)(816,1099)(935,1099){1}
//: {2}(939,1099)(951,1099){3}
//: {4}(#:937,1097)(937,1090)(1102,1090){5}
wire [31:0] w59;    //: /sn:0 {0}(#:588,629)(826,629)(826,706)(938,706){1}
//: {2}(942,706)(951,706){3}
//: {4}(#:940,704)(940,694)(978,694)(978,682)(1037,682)(1037,697)(1102,697){5}
wire w62;    //: /sn:0 {0}(8,518)(106,518)(106,394)(457,394){1}
wire w136;    //: /sn:0 {0}(-104,977)(-27,977)(-27,981)(-12,981){1}
wire w139;    //: /sn:0 {0}(-104,890)(-30,890)(-30,891)(-15,891){1}
wire w12;    //: /sn:0 {0}(6,342)(58,342)(58,128)(455,128){1}
wire [31:0] w11;    //: /sn:0 {0}(#:586,158)(912,158)(912,436)(937,436){1}
//: {2}(941,436)(951,436){3}
//: {4}(#:939,434)(939,427)(1102,427){5}
wire w137;    //: /sn:0 {0}(-104,948)(-15,948){1}
wire [31:0] w115;    //: /sn:0 {0}(#:588,1357)(833,1357)(833,1123)(933,1123){1}
//: {2}(937,1123)(951,1123){3}
//: {4}(#:935,1121)(935,1114)(1102,1114){5}
wire [31:0] w83;    //: /sn:0 {0}(#:589,1014)(687,1014)(687,927)(934,927){1}
//: {2}(938,927)(951,927){3}
//: {4}(#:936,925)(936,918)(1102,918){5}
wire w148;    //: /sn:0 {0}(-104,629)(-28,629)(-28,631)(-13,631){1}
wire w110;    //: /sn:0 {0}(457,1122)(66,1122)(66,1012)(9,1012){1}
wire w70;    //: /sn:0 {0}(458,820)(21,820)(21,807)(6,807){1}
wire w150;    //: /sn:0 {0}(-104,571)(-28,571)(-28,572)(-13,572){1}
wire [31:0] w193;    //: /sn:0 {0}(#:586,35)(932,35)(932,362)(939,362){1}
//: {2}(943,362)(#:951,362){3}
//: {4}(#:941,360)(941,353)(1102,353){5}
wire w78;    //: /sn:0 {0}(458,779)(42,779)(42,778)(6,778){1}
wire w94;    //: /sn:0 {0}(458,738)(32,738)(32,750)(6,750){1}
wire [31:0] w27;    //: /sn:0 {0}(#:586,240)(895,240)(895,485)(938,485){1}
//: {2}(942,485)(951,485){3}
//: {4}(#:940,483)(940,476)(1102,476){5}
wire [31:0] w95;    //: /sn:0 {0}(#:589,727)(811,727)(811,755)(933,755){1}
//: {2}(937,755)(951,755){3}
//: {4}(#:935,753)(935,746)(1102,746){5}
wire w86;    //: /sn:0 {0}(458,943)(95,943)(95,894)(6,894){1}
wire w138;    //: /sn:0 {0}(-104,919)(-30,919)(-30,920)(-15,920){1}
wire w142;    //: /sn:0 {0}(-104,803)(-30,803)(-30,804)(-15,804){1}
wire w155;    //: /sn:0 {0}(-104,426)(-15,426){1}
wire [31:0] w107;    //: /sn:0 {0}(#:588,1193)(735,1193)(735,1025)(932,1025){1}
//: {2}(936,1025)(951,1025){3}
//: {4}(#:934,1023)(934,1016)(1102,1016){5}
wire w143;    //: /sn:0 {0}(-104,774)(-30,774)(-30,775)(-15,775){1}
wire [31:0] w47;    //: /sn:0 {0}(#:588,424)(864,424)(864,583)(935,583){1}
//: {2}(939,583)(951,583){3}
//: {4}(#:937,581)(937,574)(1102,574){5}
wire w131;    //: /sn:0 {0}(-104,1122)(-27,1122)(-27,1125)(-12,1125){1}
wire w50;    //: /sn:0 {0}(457,681)(155,681)(155,719)(8,719){1}
wire [31:0] w79;    //: /sn:0 {0}(#:589,768)(700,768)(700,780)(932,780){1}
//: {2}(936,780)(951,780){3}
//: {4}(#:934,778)(934,771)(1102,771){5}
wire w145;    //: /sn:0 {0}(-104,716)(-13,716){1}
wire w42;    //: /sn:0 {0}(8,604)(127,604)(127,517)(457,517){1}
wire w147;    //: /sn:0 {0}(-104,658)(-28,658)(-28,659)(-13,659){1}
wire [31:0] w55;    //: /sn:0 {0}(#:588,588)(833,588)(833,681)(936,681){1}
//: {2}(940,681)(951,681){3}
//: {4}(#:938,679)(938,672)(1102,672){5}
wire [31:0] w39;    //: /sn:0 {0}(#:588,465)(855,465)(855,608)(940,608){1}
//: {2}(944,608)(951,608){3}
//: {4}(#:942,606)(942,599)(1102,599){5}
wire w26;    //: /sn:0 {0}(6,429)(83,429)(83,251)(455,251){1}
//: enddecls

  //: joint g165 (Reloj) @(413, 1277) /w:[ 8 10 -1 7 ]
  //: joint g154 (Reloj) @(413, 770) /w:[ 56 58 -1 55 ]
  Reg32bits g8 (.Din(Esc), .Reloj(Reloj), .W(w30), .Dout(w31));   //: @(456, 180) /sz:(129, 40) /sn:0 /p:[ Li0>109 Li1>109 Li2>1 Ro0<0 ]
  Decodificador5 g4 (.C(RegEsc), .S0(w160), .S1(w159), .S2(w158), .S3(w157), .S4(w156), .S5(w155), .S6(w154), .S7(w153), .S8(w152), .S9(w151), .S10(w150), .S11(w149), .S12(w148), .S13(w147), .S14(w146), .S15(w145), .S16(w144), .S17(w143), .S18(w142), .S19(w141), .S20(w140), .S21(w139), .S22(w138), .S23(w137), .S24(w136), .S25(w135), .S26(w134), .S27(w133), .S28(w132), .S29(w131), .S30(w130), .S31(w129));   //: @(-145, 252) /sz:(40, 957) /sn:0 /p:[ Li0>1 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<0 Ro6<0 Ro7<0 Ro8<0 Ro9<0 Ro10<0 Ro11<0 Ro12<0 Ro13<0 Ro14<0 Ro15<0 Ro16<0 Ro17<0 Ro18<0 Ro19<0 Ro20<0 Ro21<0 Ro22<0 Ro23<0 Ro24<0 Ro25<0 Ro26<0 Ro27<0 Ro28<0 Ro29<0 Ro30<0 Ro31<0 ]
  //: joint g186 (Esc) @(365, 800) /w:[ 52 54 -1 51 ]
  //: joint g140 (Reloj) @(413, 202) /w:[ 108 110 -1 107 ]
  Reg32bits g13 (.Din(Esc), .Reloj(Reloj), .W(w50), .Dout(w51));   //: @(458, 651) /sz:(129, 40) /sn:0 /p:[ Li0>65 Li1>65 Li2>0 Ro0<0 ]
  //: joint g37 (w15) @(940, 411) /w:[ 2 4 1 -1 ]
  //: joint g55 (w67) @(939, 853) /w:[ 1 2 4 -1 ]
  //: joint g58 (w83) @(936, 927) /w:[ 2 4 1 -1 ]
  //: joint g139 (Reloj) @(413, 161) /w:[ 112 114 -1 111 ]
  //: joint g112 (W) @(-56, 491) /w:[ 30 29 -1 32 ]
  _GGAND2 #(6) g76 (.I0(w156), .I1(W), .Z(w30));   //: @(-4,401) /sn:0 /w:[ 1 19 0 ]
  //: joint g111 (W) @(-56, 464) /w:[ 26 25 -1 28 ]
  //: joint g176 (Esc) @(365, 371) /w:[ 92 94 -1 91 ]
  //: joint g157 (Reloj) @(413, 934) /w:[ 40 42 -1 39 ]
  //: joint g163 (Reloj) @(413, 1191) /w:[ 16 18 -1 15 ]
  Reg32bits g1 (.Din(Esc), .Reloj(Reloj), .W(w4), .Dout(w7));   //: @(456, 57) /sz:(129, 40) /sn:0 /p:[ Li0>121 Li1>121 Li2>1 Ro0<0 ]
  //: joint g64 (w119) @(936, 1074) /w:[ 2 4 1 -1 ]
  //: joint g166 (Reloj) @(413, 1316) /w:[ 4 6 -1 3 ]
  Reg32bits g11 (.Din(Esc), .Reloj(Reloj), .W(w42), .Dout(w43));   //: @(458, 487) /sz:(129, 40) /sn:0 /p:[ Li0>81 Li1>81 Li2>1 Ro0<0 ]
  //: joint g130 (W) @(-56, 1022) /w:[ 102 101 -1 104 ]
  //: joint g121 (W) @(-56, 752) /w:[ 66 65 -1 68 ]
  Reg32bits g28 (.Din(Esc), .Reloj(Reloj), .W(w110), .Dout(w111));   //: @(458, 1092) /sz:(129, 40) /sn:0 /p:[ Li0>25 Li1>25 Li2>0 Ro0<0 ]
  //: joint g50 (w51) @(934, 730) /w:[ 2 4 1 -1 ]
  //: joint g197 (Esc) @(365, 1267) /w:[ 8 10 -1 7 ]
  //: joint g132 (W) @(-56, 1080) /w:[ 110 109 -1 112 ]
  Reg32bits g19 (.Din(Esc), .Reloj(Reloj), .W(w74), .Dout(w75));   //: @(459, 831) /sz:(129, 40) /sn:0 /p:[ Li0>49 Li1>49 Li2>1 Ro0<5 ]
  //: joint g113 (W) @(-56, 521) /w:[ 34 33 -1 36 ]
  //: joint g150 (Reloj) @(413, 628) /w:[ 68 70 -1 67 ]
  //: joint g146 (Reloj) @(413, 464) /w:[ 84 86 -1 83 ]
  //: joint g192 (Esc) @(365, 1060) /w:[ 28 30 -1 27 ]
  //: joint g177 (Esc) @(365, 415) /w:[ 88 90 -1 87 ]
  Reg32bits g6 (.Din(Esc), .Reloj(Reloj), .W(w22), .Dout(w23));   //: @(456, 303) /sz:(129, 40) /sn:0 /p:[ Li0>97 Li1>97 Li2>1 Ro0<0 ]
  //: joint g38 (w11) @(939, 436) /w:[ 2 4 1 -1 ]
  //: joint g115 (W) @(-56, 581) /w:[ 42 41 -1 44 ]
  Reg32bits g7 (.Din(Esc), .Reloj(Reloj), .W(w26), .Dout(w27));   //: @(456, 221) /sz:(129, 40) /sn:0 /p:[ Li0>105 Li1>105 Li2>1 Ro0<0 ]
  //: joint g53 (w71) @(936, 804) /w:[ 2 4 1 -1 ]
  _GGAND2 #(6) g75 (.I0(w157), .I1(W), .Z(w8));   //: @(-4,371) /sn:0 /w:[ 1 15 0 ]
  //: joint g169 (Esc) @(365, 67) /w:[ 120 122 -1 119 ]
  //: joint g160 (Reloj) @(413, 1073) /w:[ 28 30 -1 27 ]
  //: joint g135 (W) @(-56, 1162) /w:[ 122 121 -1 124 ]
  Reg32bits g20 (.Din(Esc), .Reloj(Reloj), .W(w78), .Dout(w79));   //: @(459, 749) /sz:(129, 40) /sn:0 /p:[ Li0>57 Li1>57 Li2>0 Ro0<0 ]
  Reg32bits g31 (.Din(Esc), .Reloj(Reloj), .W(w122), .Dout(w123));   //: @(458, 1297) /sz:(129, 40) /sn:0 /p:[ Li0>5 Li1>5 Li2>0 Ro0<0 ]
  //: joint g149 (Reloj) @(413, 589) /w:[ 72 74 -1 71 ]
  //: joint g124 (W) @(-56, 843) /w:[ 78 77 -1 80 ]
  //: joint g39 (w31) @(939, 460) /w:[ 2 4 1 -1 ]
  //: OUT g68 (Leer1) @(1263,627) /sn:0 /w:[ 0 ]
  //: joint g48 (w55) @(938, 681) /w:[ 2 4 1 -1 ]
  //: joint g195 (Esc) @(365, 1186) /w:[ 16 18 -1 15 ]
  Reg32bits g17 (.Din(Esc), .Reloj(Reloj), .W(w66), .Dout(w67));   //: @(459, 872) /sz:(129, 40) /sn:0 /p:[ Li0>45 Li1>45 Li2>0 Ro0<5 ]
  Reg32bits g25 (.Din(Esc), .Reloj(Reloj), .W(w98), .Dout(w99));   //: @(458, 1215) /sz:(129, 40) /sn:0 /p:[ Li0>13 Li1>13 Li2>1 Ro0<0 ]
  Reg32bits g29 (.Din(Esc), .Reloj(Reloj), .W(w114), .Dout(w115));   //: @(458, 1338) /sz:(129, 40) /sn:0 /p:[ Li0>0 Li1>0 Li2>0 Ro0<0 ]
  //: joint g179 (Esc) @(365, 495) /w:[ 80 82 -1 79 ]
  //: joint g52 (w79) @(934, 780) /w:[ 2 4 1 -1 ]
  //: joint g106 (W) @(-56, 313) /w:[ 6 5 -1 8 ]
  //: joint g107 (W) @(-56, 345) /w:[ 10 9 -1 12 ]
  //: joint g174 (Esc) @(365, 272) /w:[ 100 102 -1 99 ]
  _GGAND2 #(6) g83 (.I0(w146), .I1(W), .Z(w58));   //: @(-2,691) /sn:0 /w:[ 1 59 0 ]
  _GGAND2 #(6) g100 (.I0(w133), .I1(W), .Z(w106));   //: @(-1,1070) /sn:0 /w:[ 1 111 1 ]
  Reg32bits g14 (.Din(Esc), .Reloj(Reloj), .W(w54), .Dout(w55));   //: @(458, 569) /sz:(129, 40) /sn:0 /p:[ Li0>73 Li1>73 Li2>1 Ro0<0 ]
  //: joint g193 (Esc) @(365, 1102) /w:[ 24 26 -1 23 ]
  //: joint g44 (w47) @(937, 583) /w:[ 2 4 1 -1 ]
  //: joint g47 (w35) @(938, 657) /w:[ 2 4 1 -1 ]
  _GGAND2 #(6) g80 (.I0(w148), .I1(W), .Z(w34));   //: @(-2,634) /sn:0 /w:[ 1 51 0 ]
  _GGAND2 #(6) g94 (.I0(w142), .I1(W), .Z(w70));   //: @(-4,807) /sn:0 /w:[ 1 75 1 ]
  //: joint g172 (Esc) @(365, 189) /w:[ 108 110 -1 107 ]
  //: joint g159 (Reloj) @(413, 1012) /w:[ 32 34 -1 31 ]
  Reg32bits g21 (.Din(Esc), .Reloj(Reloj), .W(w82), .Dout(w83));   //: @(459, 995) /sz:(129, 40) /sn:0 /p:[ Li0>33 Li1>33 Li2>0 Ro0<0 ]
  _GGAND2 #(6) g84 (.I0(w149), .I1(W), .Z(w42));   //: @(-2,604) /sn:0 /w:[ 1 47 0 ]
  //: joint g105 (W) @(-56, 287) /w:[ 2 1 -1 4 ]
  //: joint g155 (Reloj) @(413, 850) /w:[ 48 50 -1 47 ]
  //: joint g141 (Reloj) @(413, 244) /w:[ 104 106 -1 103 ]
  Reg32bits g23 (.Din(Esc), .Reloj(Reloj), .W(w90), .Dout(w91));   //: @(459, 954) /sz:(129, 40) /sn:0 /p:[ Li0>37 Li1>37 Li2>0 Ro0<0 ]
  //: joint g41 (w19) @(936, 509) /w:[ 2 4 1 -1 ]
  //: joint g151 (Reloj) @(413, 670) /w:[ 64 66 -1 63 ]
  //: joint g40 (w27) @(940, 485) /w:[ 2 4 1 -1 ]
  //: joint g54 (w75) @(937, 829) /w:[ 1 2 4 -1 ]
  _GGAND2 #(6) g93 (.I0(w143), .I1(W), .Z(w78));   //: @(-4,778) /sn:0 /w:[ 1 71 1 ]
  //: joint g116 (W) @(-56, 612) /w:[ 46 45 -1 48 ]
  //: joint g123 (W) @(-56, 819) /w:[ 74 73 -1 76 ]
  //: joint g167 (Reloj) @(413, 1357) /w:[ 1 2 -1 124 ]
  Reg32bits g0 (.Din(Esc), .Reloj(Reloj), .W(w0), .Dout(w193));   //: @(456, 16) /sz:(129, 40) /sn:0 /p:[ Li0>123 Li1>123 Li2>1 Ro0<0 ]
  Reg32bits g26 (.Din(Esc), .Reloj(Reloj), .W(w102), .Dout(w103));   //: @(458, 1133) /sz:(129, 40) /sn:0 /p:[ Li0>21 Li1>21 Li2>0 Ro0<0 ]
  //: joint g46 (w43) @(937, 632) /w:[ 2 4 1 -1 ]
  _GGAND2 #(6) g90 (.I0(w144), .I1(W), .Z(w94));   //: @(-4,750) /sn:0 /w:[ 1 67 1 ]
  _GGAND2 #(6) g82 (.I0(w152), .I1(W), .Z(w62));   //: @(-2,518) /sn:0 /w:[ 1 35 0 ]
  //: IN g136 (Reloj) @(335,1477) /sn:0 /w:[ 125 ]
  //: joint g128 (W) @(-56, 959) /w:[ 94 93 -1 96 ]
  //: joint g190 (Esc) @(365, 967) /w:[ 36 38 -1 35 ]
  //: joint g173 (Esc) @(365, 227) /w:[ 104 106 -1 103 ]
  Mux5x32 g33 (.C(RegLeer1), .E0(w193), .E1(w7), .E2(w15), .E3(w11), .E4(w31), .E5(w27), .E6(w19), .E7(w23), .E8(w63), .E9(w47), .E10(w39), .E11(w43), .E12(w35), .E13(w55), .E14(w59), .E15(w51), .E16(w95), .E17(w79), .E18(w71), .E19(w75), .E20(w67), .E21(w87), .E22(w91), .E23(w83), .E24(w203), .E25(w111), .E26(w103), .E27(w107), .E28(w99), .E29(w119), .E30(w123), .E31(w115), .Sa(Leer1));   //: @(952, 338) /sz:(40, 835) /sn:0 /p:[ Ti0>1 Li0>3 Li1>3 Li2>3 Li3>3 Li4>3 Li5>3 Li6>3 Li7>3 Li8>3 Li9>3 Li10>3 Li11>3 Li12>3 Li13>3 Li14>3 Li15>3 Li16>3 Li17>3 Li18>3 Li19>0 Li20>0 Li21>3 Li22>3 Li23>3 Li24>3 Li25>3 Li26>3 Li27>3 Li28>3 Li29>3 Li30>3 Li31>3 Ro0<1 ]
  _GGAND2 #(6) g91 (.I0(w138), .I1(W), .Z(w90));   //: @(-4,923) /sn:0 /w:[ 1 91 1 ]
  //: joint g49 (w59) @(940, 706) /w:[ 2 4 1 -1 ]
  //: joint g198 (Esc) @(365, 1309) /w:[ 4 6 -1 3 ]
  //: joint g137 (Reloj) @(413, 75) /w:[ 120 122 -1 119 ]
  //: joint g61 (w103) @(934, 1001) /w:[ 2 4 1 -1 ]
  //: joint g158 (Reloj) @(413, 975) /w:[ 36 38 -1 35 ]
  Reg32bits g3 (.Din(Esc), .Reloj(Reloj), .W(w12), .Dout(w15));   //: @(456, 98) /sz:(129, 40) /sn:0 /p:[ Li0>117 Li1>117 Li2>1 Ro0<0 ]
  Mux5x32 g34 (.C(RegLeer2), .E0(w193), .E1(w7), .E2(w15), .E3(w11), .E4(w31), .E5(w27), .E6(w19), .E7(w23), .E8(w63), .E9(w47), .E10(w39), .E11(w43), .E12(w35), .E13(w55), .E14(w59), .E15(w51), .E16(w95), .E17(w79), .E18(w71), .E19(w75), .E20(w67), .E21(w87), .E22(w91), .E23(w83), .E24(w203), .E25(w111), .E26(w103), .E27(w107), .E28(w99), .E29(w119), .E30(w123), .E31(w115), .Sa(Leer2));   //: @(1103, 329) /sz:(40, 835) /sn:0 /p:[ Ti0>1 Li0>5 Li1>5 Li2>5 Li3>5 Li4>5 Li5>5 Li6>5 Li7>5 Li8>5 Li9>5 Li10>5 Li11>5 Li12>5 Li13>5 Li14>5 Li15>5 Li16>5 Li17>5 Li18>5 Li19>3 Li20>3 Li21>5 Li22>5 Li23>5 Li24>5 Li25>5 Li26>5 Li27>5 Li28>5 Li29>5 Li30>5 Li31>5 Ro0<0 ]
  //: joint g51 (w95) @(935, 755) /w:[ 2 4 1 -1 ]
  _GGAND2 #(6) g86 (.I0(w150), .I1(W), .Z(w38));   //: @(-2,575) /sn:0 /w:[ 1 43 0 ]
  _GGAND2 #(6) g89 (.I0(w139), .I1(W), .Z(w86));   //: @(-4,894) /sn:0 /w:[ 1 87 1 ]
  Reg32bits g2 (.Din(Esc), .Reloj(Reloj), .W(w8), .Dout(w11));   //: @(456, 139) /sz:(129, 40) /sn:0 /p:[ Li0>113 Li1>113 Li2>1 Ro0<0 ]
  //: joint g65 (w123) @(937, 1099) /w:[ 2 4 1 -1 ]
  _GGAND2 #(6) g77 (.I0(w155), .I1(W), .Z(w26));   //: @(-4,429) /sn:0 /w:[ 1 23 0 ]
  //: joint g110 (W) @(-56, 439) /w:[ 22 21 -1 24 ]
  //: joint g156 (Reloj) @(413, 892) /w:[ 44 46 -1 43 ]
  //: joint g148 (Reloj) @(413, 548) /w:[ 76 78 -1 75 ]
  //: joint g147 (Reloj) @(413, 507) /w:[ 80 82 -1 79 ]
  //: joint g59 (w203) @(937, 951) /w:[ 2 4 1 -1 ]
  //: joint g153 (Reloj) @(413, 811) /w:[ 52 54 -1 51 ]
  _GGAND2 #(6) g72 (.I0(w160), .I1(W), .Z(w0));   //: @(-4,285) /sn:0 /w:[ 1 3 0 ]
  //: joint g196 (Esc) @(365, 1227) /w:[ 12 14 -1 11 ]
  //: joint g182 (Esc) @(365, 624) /w:[ 68 70 -1 67 ]
  //: joint g161 (Reloj) @(413, 1112) /w:[ 24 26 -1 23 ]
  _GGAND2 #(6) g98 (.I0(w136), .I1(W), .Z(w126));   //: @(-1,984) /sn:0 /w:[ 1 99 1 ]
  _GGAND2 #(6) g99 (.I0(w130), .I1(W), .Z(w122));   //: @(-1,1157) /sn:0 /w:[ 1 123 1 ]
  Reg32bits g16 (.Din(Esc), .Reloj(Reloj), .W(w62), .Dout(w63));   //: @(458, 364) /sz:(129, 40) /sn:0 /p:[ Li0>93 Li1>93 Li2>1 Ro0<0 ]
  _GGAND2 #(6) g96 (.I0(w132), .I1(W), .Z(w98));   //: @(-1,1100) /sn:0 /w:[ 1 115 0 ]
  //: joint g189 (Esc) @(365, 882) /w:[ 44 46 -1 43 ]
  //: joint g183 (Esc) @(365, 718) /w:[ 60 62 -1 59 ]
  //: joint g152 (Reloj) @(413, 732) /w:[ 60 62 -1 59 ]
  _GGAND2 #(6) g103 (.I0(w129), .I1(W), .Z(w114));   //: @(-1,1185) /sn:0 /w:[ 1 125 1 ]
  //: joint g122 (W) @(-56, 786) /w:[ 70 69 -1 72 ]
  Reg32bits g10 (.Din(Esc), .Reloj(Reloj), .W(w38), .Dout(w39));   //: @(458, 446) /sz:(129, 40) /sn:0 /p:[ Li0>85 Li1>85 Li2>1 Ro0<0 ]
  _GGAND2 #(6) g78 (.I0(w154), .I1(W), .Z(w18));   //: @(-4,458) /sn:0 /w:[ 1 27 0 ]
  _GGAND2 #(6) g87 (.I0(w145), .I1(W), .Z(w50));   //: @(-2,719) /sn:0 /w:[ 1 63 1 ]
  //: joint g199 (Esc) @(365, 1353) /w:[ 1 2 -1 124 ]
  //: joint g171 (Esc) @(365, 148) /w:[ 112 114 -1 111 ]
  //: joint g129 (W) @(-56, 992) /w:[ 98 97 -1 100 ]
  Reg32bits g27 (.Din(Esc), .Reloj(Reloj), .W(w106), .Dout(w107));   //: @(458, 1174) /sz:(129, 40) /sn:0 /p:[ Li0>17 Li1>17 Li2>0 Ro0<0 ]
  Reg32bits g32 (.Din(Esc), .Reloj(Reloj), .W(w126), .Dout(w203));   //: @(458, 1051) /sz:(129, 40) /sn:0 /p:[ Li0>29 Li1>29 Li2>0 Ro0<0 ]
  //: joint g187 (Esc) @(365, 842) /w:[ 48 50 -1 47 ]
  _GGAND2 #(6) g102 (.I0(w134), .I1(W), .Z(w102));   //: @(-1,1041) /sn:0 /w:[ 1 107 1 ]
  //: joint g143 (Reloj) @(413, 323) /w:[ 96 98 -1 95 ]
  //: IN g69 (RegLeer1) @(1004,284) /sn:0 /w:[ 0 ]
  Reg32bits g9 (.Din(Esc), .Reloj(Reloj), .W(w34), .Dout(w35));   //: @(458, 528) /sz:(129, 40) /sn:0 /p:[ Li0>77 Li1>77 Li2>1 Ro0<0 ]
  //: joint g57 (w91) @(937, 902) /w:[ 2 4 1 -1 ]
  //: joint g119 (W) @(-56, 698) /w:[ 58 57 -1 60 ]
  //: joint g142 (Reloj) @(413, 282) /w:[ 100 102 -1 99 ]
  Reg32bits g15 (.Din(Esc), .Reloj(Reloj), .W(w58), .Dout(w59));   //: @(458, 610) /sz:(129, 40) /sn:0 /p:[ Li0>69 Li1>69 Li2>1 Ro0<0 ]
  //: IN g71 (RegEsc) @(-281,700) /sn:0 /w:[ 0 ]
  //: joint g162 (Reloj) @(413, 1153) /w:[ 20 22 -1 19 ]
  //: joint g131 (W) @(-56, 1047) /w:[ 106 105 -1 108 ]
  //: OUT g67 (Leer2) @(1263,687) /sn:0 /w:[ 1 ]
  //: joint g127 (W) @(-56, 930) /w:[ 90 89 -1 92 ]
  //: joint g43 (w63) @(937, 559) /w:[ 2 4 1 -1 ]
  //: joint g145 (Reloj) @(413, 423) /w:[ 88 90 -1 87 ]
  //: joint g62 (w107) @(934, 1025) /w:[ 2 4 1 -1 ]
  _GGAND2 #(6) g73 (.I0(w159), .I1(W), .Z(w4));   //: @(-4,313) /sn:0 /w:[ 1 7 0 ]
  _GGAND2 #(6) g88 (.I0(w140), .I1(W), .Z(w66));   //: @(-4,866) /sn:0 /w:[ 1 83 1 ]
  //: IN g104 (W) @(-143,203) /sn:0 /w:[ 0 ]
  //: joint g188 (Esc) @(365, 922) /w:[ 40 42 -1 39 ]
  //: joint g180 (Esc) @(365, 536) /w:[ 76 78 -1 75 ]
  //: joint g138 (Reloj) @(413, 116) /w:[ 116 118 -1 115 ]
  //: joint g42 (w23) @(935, 534) /w:[ 2 4 1 -1 ]
  //: joint g63 (w99) @(937, 1050) /w:[ 2 4 1 -1 ]
  //: joint g175 (Esc) @(365, 311) /w:[ 96 98 -1 95 ]
  _GGAND2 #(6) g74 (.I0(w158), .I1(W), .Z(w12));   //: @(-4,342) /sn:0 /w:[ 1 11 0 ]
  //: joint g109 (W) @(-56, 410) /w:[ 18 17 -1 20 ]
  //: joint g181 (Esc) @(365, 579) /w:[ 72 74 -1 71 ]
  //: IN g168 (Esc) @(324,1422) /sn:0 /w:[ 125 ]
  //: joint g133 (W) @(-56, 1105) /w:[ 114 113 -1 116 ]
  Reg32bits g5 (.Din(Esc), .Reloj(Reloj), .W(w18), .Dout(w19));   //: @(456, 262) /sz:(129, 40) /sn:0 /p:[ Li0>101 Li1>101 Li2>1 Ro0<0 ]
  //: joint g56 (w87) @(936, 878) /w:[ 2 4 1 -1 ]
  //: joint g194 (Esc) @(365, 1143) /w:[ 20 22 -1 19 ]
  _GGAND2 #(6) g79 (.I0(w153), .I1(W), .Z(w22));   //: @(-4,486) /sn:0 /w:[ 1 31 0 ]
  _GGAND2 #(6) g95 (.I0(w137), .I1(W), .Z(w82));   //: @(-4,951) /sn:0 /w:[ 1 95 1 ]
  //: joint g117 (W) @(-56, 640) /w:[ 50 49 -1 52 ]
  Reg32bits g24 (.Din(Esc), .Reloj(Reloj), .W(w94), .Dout(w95));   //: @(459, 708) /sz:(129, 40) /sn:0 /p:[ Li0>61 Li1>61 Li2>0 Ro0<0 ]
  //: joint g36 (w7) @(939, 387) /w:[ 2 4 1 -1 ]
  _GGAND2 #(6) g85 (.I0(w151), .I1(W), .Z(w46));   //: @(-2,546) /sn:0 /w:[ 1 39 0 ]
  _GGAND2 #(6) g92 (.I0(w141), .I1(W), .Z(w74));   //: @(-4,836) /sn:0 /w:[ 1 79 0 ]
  //: joint g178 (Esc) @(365, 455) /w:[ 84 86 -1 83 ]
  //: joint g144 (Reloj) @(413, 384) /w:[ 92 94 -1 91 ]
  //: joint g125 (W) @(-56, 874) /w:[ 82 81 -1 84 ]
  //: joint g60 (w111) @(935, 976) /w:[ 2 4 1 -1 ]
  _GGAND2 #(6) g81 (.I0(w147), .I1(W), .Z(w54));   //: @(-2,662) /sn:0 /w:[ 1 55 0 ]
  _GGAND2 #(6) g101 (.I0(w135), .I1(W), .Z(w110));   //: @(-1,1012) /sn:0 /w:[ 1 103 1 ]
  //: joint g185 (Esc) @(365, 763) /w:[ 56 58 -1 55 ]
  //: joint g170 (Esc) @(365, 107) /w:[ 116 118 -1 115 ]
  Reg32bits g22 (.Din(Esc), .Reloj(Reloj), .W(w86), .Dout(w87));   //: @(459, 913) /sz:(129, 40) /sn:0 /p:[ Li0>41 Li1>41 Li2>0 Ro0<0 ]
  //: joint g35 (w193) @(941, 362) /w:[ 2 4 1 -1 ]
  //: joint g45 (w39) @(942, 608) /w:[ 2 4 1 -1 ]
  //: IN g70 (RegLeer2) @(1145,282) /sn:0 /w:[ 0 ]
  //: joint g126 (W) @(-56, 903) /w:[ 86 85 -1 88 ]
  //: joint g184 (Esc) @(365, 661) /w:[ 64 66 -1 63 ]
  //: joint g66 (w115) @(935, 1123) /w:[ 2 4 1 -1 ]
  _GGAND2 #(6) g97 (.I0(w131), .I1(W), .Z(w118));   //: @(-1,1128) /sn:0 /w:[ 1 119 1 ]
  //: joint g114 (W) @(-56, 553) /w:[ 38 37 -1 40 ]
  //: joint g120 (W) @(-56, 725) /w:[ 62 61 -1 64 ]
  Reg32bits g12 (.Din(Esc), .Reloj(Reloj), .W(w46), .Dout(w47));   //: @(458, 405) /sz:(129, 40) /sn:0 /p:[ Li0>89 Li1>89 Li2>1 Ro0<0 ]
  Reg32bits g18 (.Din(Esc), .Reloj(Reloj), .W(w70), .Dout(w71));   //: @(459, 790) /sz:(129, 40) /sn:0 /p:[ Li0>53 Li1>53 Li2>0 Ro0<0 ]
  //: joint g191 (Esc) @(365, 1005) /w:[ 32 34 -1 31 ]
  //: joint g164 (Reloj) @(413, 1235) /w:[ 12 14 -1 11 ]
  Reg32bits g30 (.Din(Esc), .Reloj(Reloj), .W(w118), .Dout(w119));   //: @(458, 1256) /sz:(129, 40) /sn:0 /p:[ Li0>9 Li1>9 Li2>0 Ro0<0 ]
  //: joint g108 (W) @(-56, 377) /w:[ 14 13 -1 16 ]
  //: joint g134 (W) @(-56, 1134) /w:[ 118 117 -1 120 ]
  //: joint g118 (W) @(-56, 669) /w:[ 54 53 -1 56 ]

endmodule
//: /netlistEnd

//: /netlistBegin Reg32bits
module Reg32bits(W, Reloj, Dout, Din);
//: interface  /sz:(97, 40) /bd:[ Li0>W(30/40) Li1>Reloj(20/40) Li2>Din[31:0](10/40) Ro0<Dout[31:0](19/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [31:0] Din;    //: /sn:0 {0}(#:12,40)(54,40)(54,41)(#:69,41){1}
output [31:0] Dout;    //: /sn:0 {0}(#:3199,423)(3323,423){1}
input Reloj;    //: /sn:0 {0}(2833,220)(2824,220)(2824,282){1}
//: {2}(2826,284)(2908,284){3}
//: {4}(2912,284)(2990,284){5}
//: {6}(2994,284)(3080,284)(3080,220)(3095,220){7}
//: {8}(2992,282)(2992,221)(3006,221){9}
//: {10}(2910,282)(2910,222)(2921,222){11}
//: {12}(2822,284)(2736,284){13}
//: {14}(2734,282)(2734,221)(2747,221){15}
//: {16}(2732,284)(2646,284){17}
//: {18}(2644,282)(2644,222)(2658,222){19}
//: {20}(2642,284)(2564,284){21}
//: {22}(2562,282)(2562,223)(2573,223){23}
//: {24}(2560,284)(2473,284){25}
//: {26}(2471,282)(2471,221)(2485,221){27}
//: {28}(2469,284)(2307,284){29}
//: {30}(2305,282)(2305,222)(2319,222){31}
//: {32}(2303,284)(2210,284){33}
//: {34}(2208,282)(2208,223)(2230,223){35}
//: {36}(2206,284)(2131,284){37}
//: {38}(2129,282)(2129,224)(2145,224){39}
//: {40}(2127,284)(2046,284){41}
//: {42}(2044,282)(2044,222)(2057,222){43}
//: {44}(2042,284)(1960,284){45}
//: {46}(1958,282)(1958,223)(1971,223){47}
//: {48}(1956,284)(1878,284){49}
//: {50}(1876,282)(1876,224)(1882,224){51}
//: {52}(1874,284)(1788,284){53}
//: {54}(1786,282)(1786,225)(1797,225){55}
//: {56}(1784,284)(1692,284){57}
//: {58}(1690,282)(1690,223)(1709,223){59}
//: {60}(1688,284)(1536,284){61}
//: {62}(1534,282)(1534,225)(1541,225){63}
//: {64}(1532,284)(1444,284){65}
//: {66}(1442,282)(1442,226)(1452,226){67}
//: {68}(1440,284)(1354,284){69}
//: {70}(1352,282)(1352,227)(1367,227){71}
//: {72}(1350,284)(1268,284){73}
//: {74}(1266,282)(1266,225)(1279,225){75}
//: {76}(1264,284)(1186,284){77}
//: {78}(1184,282)(1184,226)(1193,226){79}
//: {80}(1182,284)(1097,284){81}
//: {82}(1095,282)(1095,227)(1104,227){83}
//: {84}(1093,284)(1010,284){85}
//: {86}(1008,282)(1008,228)(1019,228){87}
//: {88}(1006,284)(922,284){89}
//: {90}(920,282)(920,226)(931,226){91}
//: {92}(918,284)(733,284){93}
//: {94}(731,282)(731,226)(741,226){95}
//: {96}(729,284)(643,284){97}
//: {98}(641,282)(641,227)(652,227){99}
//: {100}(639,284)(554,284){101}
//: {102}(552,282)(552,228)(567,228){103}
//: {104}(550,284)(468,284){105}
//: {106}(466,282)(466,226)(479,226){107}
//: {108}(464,284)(387,284){109}
//: {110}(385,282)(385,227)(393,227){111}
//: {112}(383,284)(294,284){113}
//: {114}(292,282)(292,228)(304,228){115}
//: {116}(290,284)(211,284){117}
//: {118}(209,282)(209,229)(219,229){119}
//: {120}(207,284)(118,284){121}
//: {122}(116,282)(116,227)(131,227){123}
//: {124}(114,284)(2,284){125}
input W;    //: /sn:0 {0}(3040,233)(3040,302)(3037,302)(3037,312){1}
//: {2}(3039,314)(3129,314)(3129,232){3}
//: {4}(3035,314)(2958,314){5}
//: {6}(2956,312)(2956,302)(2955,302)(2955,234){7}
//: {8}(2954,314)(2867,314){9}
//: {10}(2865,312)(2865,302)(2867,302)(2867,232){11}
//: {12}(2863,314)(2781,314){13}
//: {14}(2779,312)(2779,302)(2781,302)(2781,233){15}
//: {16}(2777,314)(2695,314){17}
//: {18}(2693,312)(2693,302)(2692,302)(2692,234){19}
//: {20}(2691,314)(2608,314){21}
//: {22}(2606,312)(2606,302)(2607,302)(2607,235){23}
//: {24}(2604,314)(2519,314){25}
//: {26}(2517,312)(2517,302)(2519,302)(2519,233){27}
//: {28}(2515,314)(2355,314){29}
//: {30}(2353,312)(2353,234){31}
//: {32}(2351,314)(2267,314){33}
//: {34}(2265,312)(2265,302)(2264,302)(2264,235){35}
//: {36}(2263,314)(2173,314){37}
//: {38}(2171,312)(2171,302)(2179,302)(2179,236){39}
//: {40}(2169,314)(2090,314){41}
//: {42}(2088,312)(2088,302)(2091,302)(2091,234){43}
//: {44}(2086,314)(2007,314){45}
//: {46}(2005,312)(2005,235){47}
//: {48}(2003,314)(1918,314){49}
//: {50}(1916,312)(1916,236){51}
//: {52}(1914,314)(1827,314){53}
//: {54}(1825,312)(1825,302)(1831,302)(1831,237){55}
//: {56}(1823,314)(1737,314){57}
//: {58}(1735,312)(1735,302)(1743,302)(1743,235){59}
//: {60}(1733,314)(1576,314){61}
//: {62}(1574,312)(1574,302)(1575,302)(1575,237){63}
//: {64}(1572,314)(1484,314){65}
//: {66}(1482,312)(1482,302)(1486,302)(1486,238){67}
//: {68}(1480,314)(1404,314){69}
//: {70}(1402,312)(1402,302)(1401,302)(1401,239){71}
//: {72}(1400,314)(1314,314){73}
//: {74}(1312,312)(1312,302)(1313,302)(1313,237){75}
//: {76}(1310,314)(1229,314){77}
//: {78}(1227,312)(1227,238){79}
//: {80}(1225,314)(1142,314){81}
//: {82}(1140,312)(1140,302)(1138,302)(1138,239){83}
//: {84}(1138,314)(1057,314){85}
//: {86}(1055,312)(1055,302)(1053,302)(1053,240){87}
//: {88}(1053,314)(964,314){89}
//: {90}(962,312)(962,302)(965,302)(965,238){91}
//: {92}(960,314)(774,314){93}
//: {94}(772,312)(772,302)(775,302)(775,238){95}
//: {96}(770,314)(688,314){97}
//: {98}(686,312)(686,239){99}
//: {100}(684,314)(607,314){101}
//: {102}(605,312)(605,302)(601,302)(601,240){103}
//: {104}(603,314)(517,314){105}
//: {106}(515,312)(515,302)(513,302)(513,238){107}
//: {108}(513,314)(430,314){109}
//: {110}(428,312)(428,302)(427,302)(427,239){111}
//: {112}(426,314)(340,314){113}
//: {114}(338,312)(338,240){115}
//: {116}(336,314)(257,314){117}
//: {118}(255,312)(255,302)(253,302)(253,241){119}
//: {120}(253,314)(170,314){121}
//: {122}(168,312)(168,302)(165,302)(165,239){123}
//: {124}(166,314)(0,314){125}
wire w73;    //: /sn:0 {0}(1321,215)(1336,215){1}
wire w96;    //: /sn:0 {0}(2230,200)(2214,200)(2214,115)(2074,115)(2074,91){1}
wire w93;    //: /sn:0 {0}(1751,213)(1766,213){1}
wire w134;    //: /sn:0 {0}(2527,197)(2550,197)(2550,352)(2822,352)(2822,375){1}
wire w46;    //: /sn:0 {0}(1367,204)(1348,204)(1348,127)(1296,127)(1296,95){1}
wire w61;    //: /sn:0 {0}(1316,95)(1316,113)(1524,113)(1524,202)(1541,202){1}
wire w99;    //: /sn:0 {0}(2272,199)(2294,199)(2294,347)(2134,347)(2134,376){1}
wire w141;    //: /sn:0 {0}(2867,96)(2867,116)(3081,116)(3081,197)(3095,197){1}
wire w14;    //: /sn:0 {0}(346,218)(361,218){1}
wire w56;    //: /sn:0 {0}(1452,203)(1433,203)(1433,120)(1306,120)(1306,95){1}
wire w153;    //: /sn:0 {0}(2875,210)(2890,210){1}
wire w4;    //: /sn:0 {0}(173,217)(188,217){1}
wire w19;    //: /sn:0 {0}(435,217)(450,217){1}
wire w81;    //: /sn:0 {0}(1797,202)(1787,202)(1787,134)(2024,134)(2024,91){1}
wire w89;    //: /sn:0 {0}(2187,200)(2197,200)(2197,341)(2124,341)(2124,376){1}
wire w15;    //: /sn:0 {0}(393,204)(383,204)(383,174)(469,174)(469,125){1}
wire [7:0] w195;    //: /sn:0 {0}(#:75,56)(474,56)(#:474,119){1}
wire w38;    //: /sn:0 {0}(694,217)(709,217){1}
wire [7:0] w213;    //: /sn:0 {0}(3193,428)(2109,428)(#:2109,382){1}
wire w129;    //: /sn:0 {0}(2963,198)(2983,198)(2983,337)(2872,337)(2872,375){1}
wire w51;    //: /sn:0 {0}(931,203)(921,203)(921,123)(1246,123)(1246,95){1}
wire w69;    //: /sn:0 {0}(1292,396)(1292,350)(1258,350)(1258,202)(1235,202){1}
wire w106;    //: /sn:0 {0}(1971,200)(1955,200)(1955,152)(2044,152)(2044,91){1}
wire w109;    //: /sn:0 {0}(2104,376)(2104,335)(2035,335)(2035,199)(2013,199){1}
wire w151;    //: /sn:0 {0}(2833,197)(2821,197)(2821,181)(2837,181)(2837,96){1}
wire w0;    //: /sn:0 {0}(131,204)(121,204)(121,160)(439,160)(439,125){1}
wire w3;    //: /sn:0 {0}(445,382)(445,353)(197,353)(197,203)(173,203){1}
wire w114;    //: /sn:0 {0}(2114,376)(2114,337)(2121,337)(2121,198)(2099,198){1}
wire w128;    //: /sn:0 {0}(2963,212)(2978,212){1}
wire [7:0] w177;    //: /sn:0 {0}(75,36)(2049,36)(#:2049,85){1}
wire w64;    //: /sn:0 {0}(1332,396)(1332,373)(1606,373)(1606,201)(1583,201){1}
wire w66;    //: /sn:0 {0}(1193,203)(1178,203)(1178,143)(1276,143)(1276,95){1}
wire w133;    //: /sn:0 {0}(2527,211)(2542,211){1}
wire w104;    //: /sn:0 {0}(2361,198)(2421,198)(2421,356)(2144,356)(2144,376){1}
wire w111;    //: /sn:0 {0}(2057,199)(2040,199)(2040,163)(2054,163)(2054,91){1}
wire w159;    //: /sn:0 {0}(2842,375)(2842,331)(2728,331)(2728,198)(2700,198){1}
wire w34;    //: /sn:0 {0}(515,382)(515,360)(809,360)(809,202)(783,202){1}
wire w63;    //: /sn:0 {0}(1583,215)(1598,215){1}
wire [7:0] w204;    //: /sn:0 {0}(3193,438)(2857,438)(#:2857,381){1}
wire w21;    //: /sn:0 {0}(489,125)(489,157)(549,157)(549,205)(567,205){1}
wire w43;    //: /sn:0 {0}(1061,218)(1076,218){1}
wire w76;    //: /sn:0 {0}(1104,204)(1094,204)(1094,134)(1266,134)(1266,95){1}
wire w54;    //: /sn:0 {0}(1262,396)(1262,368)(992,368)(992,202)(973,202){1}
wire w119;    //: /sn:0 {0}(2094,376)(2094,339)(1950,339)(1950,200)(1924,200){1}
wire w31;    //: /sn:0 {0}(509,125)(509,143)(719,143)(719,203)(741,203){1}
wire w58;    //: /sn:0 {0}(1494,216)(1509,216){1}
wire w156;    //: /sn:0 {0}(2658,199)(2648,199)(2648,162)(2817,162)(2817,96){1}
wire w28;    //: /sn:0 {0}(521,216)(536,216){1}
wire w23;    //: /sn:0 {0}(609,218)(624,218){1}
wire w36;    //: /sn:0 {0}(499,125)(499,150)(640,150)(640,204)(652,204){1}
wire w41;    //: /sn:0 {0}(1019,205)(1009,205)(1009,127)(1256,127)(1256,95){1}
wire w124;    //: /sn:0 {0}(2615,199)(2637,199)(2637,341)(2832,341)(2832,375){1}
wire w24;    //: /sn:0 {0}(495,382)(495,345)(630,345)(630,204)(609,204){1}
wire w108;    //: /sn:0 {0}(2013,213)(2028,213){1}
wire w126;    //: /sn:0 {0}(2921,199)(2906,199)(2906,135)(2847,135)(2847,96){1}
wire w154;    //: /sn:0 {0}(2862,375)(2862,325)(2898,325)(2898,196)(2875,196){1}
wire w158;    //: /sn:0 {0}(2700,212)(2715,212){1}
wire w74;    //: /sn:0 {0}(1302,396)(1302,349)(1341,349)(1341,201)(1321,201){1}
wire w98;    //: /sn:0 {0}(2272,213)(2287,213){1}
wire w116;    //: /sn:0 {0}(1882,201)(1867,201)(1867,142)(2034,142)(2034,91){1}
wire w8;    //: /sn:0 {0}(455,382)(455,348)(284,348)(284,205)(261,205){1}
wire w91;    //: /sn:0 {0}(1709,200)(1699,200)(1699,125)(2014,125)(2014,91){1}
wire w103;    //: /sn:0 {0}(2361,212)(2376,212){1}
wire w18;    //: /sn:0 {0}(475,382)(475,339)(455,339)(455,203)(435,203){1}
wire w118;    //: /sn:0 {0}(1924,214)(1939,214){1}
wire w121;    //: /sn:0 {0}(2573,200)(2563,200)(2563,150)(2807,150)(2807,96){1}
wire w71;    //: /sn:0 {0}(1279,202)(1269,202)(1269,148)(1286,148)(1286,95){1}
wire w101;    //: /sn:0 {0}(2084,91)(2084,107)(2302,107)(2302,199)(2319,199){1}
wire [7:0] w162;    //: /sn:0 {0}(75,26)(2832,26)(#:2832,90){1}
wire w68;    //: /sn:0 {0}(1235,216)(1250,216){1}
wire w144;    //: /sn:0 {0}(3137,196)(3169,196)(3169,355)(2892,355)(2892,375){1}
wire [7:0] w222;    //: /sn:0 {0}(#:3193,418)(1297,418)(#:1297,402){1}
wire w149;    //: /sn:0 {0}(2789,197)(2816,197)(2816,323)(2852,323)(2852,375){1}
wire w146;    //: /sn:0 {0}(2747,198)(2736,198)(2736,172)(2827,172)(2827,96){1}
wire w53;    //: /sn:0 {0}(973,216)(988,216){1}
wire w84;    //: /sn:0 {0}(2084,376)(2084,345)(1862,345)(1862,201)(1839,201){1}
wire w59;    //: /sn:0 {0}(1322,396)(1322,364)(1515,364)(1515,202)(1494,202){1}
wire w123;    //: /sn:0 {0}(2615,213)(2630,213){1}
wire w44;    //: /sn:0 {0}(1272,396)(1272,359)(1085,359)(1085,204)(1061,204){1}
wire w113;    //: /sn:0 {0}(2099,212)(2114,212){1}
wire w197;    //: /sn:0 {0}(2882,375)(2882,346)(3071,346)(3071,197)(3048,197){1}
wire w136;    //: /sn:0 {0}(3006,198)(2993,198)(2993,126)(2857,126)(2857,96){1}
wire w49;    //: /sn:0 {0}(1312,396)(1312,358)(1428,358)(1428,203)(1409,203){1}
wire w83;    //: /sn:0 {0}(1839,215)(1854,215){1}
wire w148;    //: /sn:0 {0}(2789,211)(2804,211){1}
wire w10;    //: /sn:0 {0}(304,205)(294,205)(294,171)(459,171)(459,125){1}
wire w78;    //: /sn:0 {0}(1146,217)(1161,217){1}
wire [7:0] w186;    //: /sn:0 {0}(#:75,46)(1281,46)(#:1281,89){1}
wire w13;    //: /sn:0 {0}(465,382)(465,344)(373,344)(373,204)(346,204){1}
wire w88;    //: /sn:0 {0}(2187,214)(2202,214){1}
wire w94;    //: /sn:0 {0}(2074,376)(2074,351)(1776,351)(1776,199)(1751,199){1}
wire w138;    //: /sn:0 {0}(3048,211)(3063,211){1}
wire w86;    //: /sn:0 {0}(2064,91)(2064,122)(2127,122)(2127,201)(2145,201){1}
wire w5;    //: /sn:0 {0}(219,206)(209,206)(209,166)(449,166)(449,125){1}
wire w33;    //: /sn:0 {0}(783,216)(798,216){1}
wire w48;    //: /sn:0 {0}(1409,217)(1424,217){1}
wire [7:0] w231;    //: /sn:0 {0}(#:3193,408)(480,408)(#:480,388){1}
wire w29;    //: /sn:0 {0}(485,382)(485,340)(543,340)(543,202)(521,202){1}
wire w143;    //: /sn:0 {0}(3137,210)(3152,210){1}
wire w131;    //: /sn:0 {0}(2485,198)(2475,198)(2475,137)(2797,137)(2797,96){1}
wire w9;    //: /sn:0 {0}(261,219)(276,219){1}
wire w79;    //: /sn:0 {0}(1282,396)(1282,355)(1170,355)(1170,203)(1146,203){1}
wire w26;    //: /sn:0 {0}(479,125)(479,180)(469,180)(469,203)(479,203){1}
wire w39;    //: /sn:0 {0}(694,203)(715,203)(715,351)(505,351)(505,382){1}
//: enddecls

  //: joint g61 (Reloj) @(1442, 284) /w:[ 65 66 68 -1 ]
  FlipFlopD g8 (.Reloj(Reloj), .D(w21), .W(W), .nQ(w23), .Q(w24));   //: @(568, 199) /sz:(40, 40) /sn:0 /p:[ Li0>103 Li1>1 Bi0>103 Ro0<0 Ro1<1 ]
  FlipFlopD g4 (.Reloj(Reloj), .D(w5), .W(W), .nQ(w9), .Q(w8));   //: @(220, 200) /sz:(40, 40) /sn:0 /p:[ Li0>119 Li1>0 Bi0>119 Ro0<0 Ro1<1 ]
  //: joint g86 (W) @(1055, 314) /w:[ 85 86 88 -1 ]
  //: joint g58 (Reloj) @(1184, 284) /w:[ 77 78 80 -1 ]
  //: joint g55 (Reloj) @(920, 284) /w:[ 89 90 92 -1 ]
  //: joint g51 (Reloj) @(466, 284) /w:[ 105 106 108 -1 ]
  assign {w91, w81, w116, w106, w111, w86, w96, w101} = w177; //: CONCAT g37  @(2049,86) /sn:0 /R:1 /w:[ 1 1 1 1 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  FlipFlopD g34 (.Reloj(Reloj), .D(w151), .W(W), .nQ(w153), .Q(w154));   //: @(2834, 191) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>0 Bi0>11 Ro0<0 Ro1<1 ]
  FlipFlopD g13 (.Reloj(Reloj), .D(w46), .W(W), .nQ(w48), .Q(w49));   //: @(1368, 198) /sz:(40, 40) /sn:0 /p:[ Li0>71 Li1>0 Bi0>71 Ro0<0 Ro1<1 ]
  FlipFlopD g3 (.Reloj(Reloj), .D(w0), .W(W), .nQ(w4), .Q(w3));   //: @(132, 198) /sz:(40, 40) /sn:0 /p:[ Li0>123 Li1>0 Bi0>123 Ro0<0 Ro1<1 ]
  //: joint g89 (W) @(1312, 314) /w:[ 73 74 76 -1 ]
  //: joint g77 (W) @(168, 314) /w:[ 121 122 124 -1 ]
  //: joint g76 (Reloj) @(2910, 284) /w:[ 4 10 3 -1 ]
  //: joint g65 (Reloj) @(1876, 284) /w:[ 49 50 52 -1 ]
  //: IN g2 (W) @(-2,314) /sn:0 /w:[ 125 ]
  //: joint g59 (Reloj) @(1266, 284) /w:[ 73 74 76 -1 ]
  //: joint g72 (Reloj) @(2562, 284) /w:[ 21 22 24 -1 ]
  //: IN g1 (Reloj) @(0,284) /sn:0 /w:[ 125 ]
  //: joint g99 (W) @(2265, 314) /w:[ 33 34 36 -1 ]
  //: joint g98 (W) @(2171, 314) /w:[ 37 38 40 -1 ]
  //: joint g64 (Reloj) @(1786, 284) /w:[ 53 54 56 -1 ]
  //: joint g96 (W) @(2005, 314) /w:[ 45 46 48 -1 ]
  FlipFlopD g16 (.Reloj(Reloj), .D(w61), .W(W), .nQ(w63), .Q(w64));   //: @(1542, 196) /sz:(40, 40) /sn:0 /p:[ Li0>63 Li1>1 Bi0>63 Ro0<0 Ro1<1 ]
  FlipFlopD g11 (.Reloj(Reloj), .D(w36), .W(W), .nQ(w38), .Q(w39));   //: @(653, 198) /sz:(40, 40) /sn:0 /p:[ Li0>99 Li1>1 Bi0>99 Ro0<0 Ro1<0 ]
  //: joint g103 (W) @(2693, 314) /w:[ 17 18 20 -1 ]
  //: joint g87 (W) @(1140, 314) /w:[ 81 82 84 -1 ]
  //: joint g78 (W) @(255, 314) /w:[ 117 118 120 -1 ]
  //: joint g50 (Reloj) @(385, 284) /w:[ 109 110 112 -1 ]
  FlipFlopD g28 (.Reloj(Reloj), .D(w121), .W(W), .nQ(w123), .Q(w124));   //: @(2574, 194) /sz:(40, 40) /sn:0 /p:[ Li0>23 Li1>0 Bi0>23 Ro0<0 Ro1<0 ]
  FlipFlopD g10 (.Reloj(Reloj), .D(w31), .W(W), .nQ(w33), .Q(w34));   //: @(742, 197) /sz:(40, 40) /sn:0 /p:[ Li0>95 Li1>1 Bi0>95 Ro0<0 Ro1<1 ]
  FlipFlopD g32 (.Reloj(Reloj), .D(w141), .W(W), .nQ(w143), .Q(w144));   //: @(3096, 191) /sz:(40, 40) /sn:0 /p:[ Li0>7 Li1>1 Bi0>3 Ro0<0 Ro1<0 ]
  FlipFlopD g27 (.Reloj(Reloj), .D(w116), .W(W), .nQ(w118), .Q(w119));   //: @(1883, 195) /sz:(40, 40) /sn:0 /p:[ Li0>51 Li1>0 Bi0>51 Ro0<0 Ro1<1 ]
  FlipFlopD g19 (.Reloj(Reloj), .D(w76), .W(W), .nQ(w78), .Q(w79));   //: @(1105, 198) /sz:(40, 40) /sn:0 /p:[ Li0>83 Li1>0 Bi0>83 Ro0<0 Ro1<1 ]
  //: joint g102 (W) @(2606, 314) /w:[ 21 22 24 -1 ]
  //: joint g69 (Reloj) @(2208, 284) /w:[ 33 34 36 -1 ]
  assign {w51, w41, w76, w66, w71, w46, w56, w61} = w186; //: CONCAT g38  @(1281,90) /sn:0 /R:1 /w:[ 1 1 1 1 1 1 1 0 1 ] /dr:0 /tp:0 /drp:0
  FlipFlopD g6 (.Reloj(Reloj), .D(w15), .W(W), .nQ(w19), .Q(w18));   //: @(394, 198) /sz:(40, 40) /sn:0 /p:[ Li0>111 Li1>0 Bi0>111 Ro0<0 Ro1<1 ]
  //: joint g75 (Reloj) @(2824, 284) /w:[ 2 1 12 -1 ]
  //: joint g57 (Reloj) @(1095, 284) /w:[ 81 82 84 -1 ]
  //: joint g53 (Reloj) @(641, 284) /w:[ 97 98 100 -1 ]
  //: OUT g7 (Dout) @(3320,423) /sn:0 /w:[ 1 ]
  FlipFlopD g9 (.Reloj(Reloj), .D(w26), .W(W), .nQ(w28), .Q(w29));   //: @(480, 197) /sz:(40, 40) /sn:0 /p:[ Li0>107 Li1>1 Bi0>107 Ro0<0 Ro1<1 ]
  //: joint g71 (Reloj) @(2471, 284) /w:[ 25 26 28 -1 ]
  FlipFlopD g31 (.Reloj(Reloj), .D(w136), .W(W), .nQ(w138), .Q(w197));   //: @(3007, 192) /sz:(40, 40) /sn:0 /p:[ Li0>9 Li1>0 Bi0>0 Ro0<0 Ro1<1 ]
  FlipFlopD g20 (.Reloj(Reloj), .D(w81), .W(W), .nQ(w83), .Q(w84));   //: @(1798, 196) /sz:(40, 40) /sn:0 /p:[ Li0>55 Li1>0 Bi0>55 Ro0<0 Ro1<1 ]
  FlipFlopD g15 (.Reloj(Reloj), .D(w56), .W(W), .nQ(w58), .Q(w59));   //: @(1453, 197) /sz:(40, 40) /sn:0 /p:[ Li0>67 Li1>0 Bi0>67 Ro0<0 Ro1<1 ]
  //: joint g68 (Reloj) @(2129, 284) /w:[ 37 38 40 -1 ]
  //: joint g67 (Reloj) @(2044, 284) /w:[ 41 42 44 -1 ]
  assign {w0, w5, w10, w15, w26, w21, w36, w31} = w195; //: CONCAT g39  @(474,120) /sn:0 /R:1 /w:[ 1 1 1 1 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: joint g48 (Reloj) @(209, 284) /w:[ 117 118 120 -1 ]
  assign w231 = {w3, w8, w13, w18, w29, w24, w39, w34}; //: CONCAT g43  @(480,387) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 1 0 ] /dr:1 /tp:0 /drp:1
  //: joint g104 (W) @(2779, 314) /w:[ 13 14 16 -1 ]
  //: joint g88 (W) @(1227, 314) /w:[ 77 78 80 -1 ]
  //: joint g73 (Reloj) @(2644, 284) /w:[ 17 18 20 -1 ]
  //: joint g62 (Reloj) @(1534, 284) /w:[ 61 62 64 -1 ]
  FlipFlopD g29 (.Reloj(Reloj), .D(w126), .W(W), .nQ(w128), .Q(w129));   //: @(2922, 193) /sz:(40, 40) /sn:0 /p:[ Li0>11 Li1>0 Bi0>7 Ro0<0 Ro1<0 ]
  FlipFlopD g25 (.Reloj(Reloj), .D(w106), .W(W), .nQ(w108), .Q(w109));   //: @(1972, 194) /sz:(40, 40) /sn:0 /p:[ Li0>47 Li1>0 Bi0>47 Ro0<0 Ro1<1 ]
  FlipFlopD g17 (.Reloj(Reloj), .D(w66), .W(W), .nQ(w68), .Q(w69));   //: @(1194, 197) /sz:(40, 40) /sn:0 /p:[ Li0>79 Li1>0 Bi0>79 Ro0<0 Ro1<1 ]
  //: joint g107 (W) @(3037, 314) /w:[ 2 1 4 -1 ]
  //: joint g106 (W) @(2956, 314) /w:[ 5 6 8 -1 ]
  //: joint g63 (Reloj) @(1690, 284) /w:[ 57 58 60 -1 ]
  //: joint g52 (Reloj) @(552, 284) /w:[ 101 102 104 -1 ]
  assign w222 = {w54, w44, w79, w69, w74, w49, w59, w64}; //: CONCAT g42  @(1297,401) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 0 0 ] /dr:1 /tp:0 /drp:1
  //: joint g83 (W) @(686, 314) /w:[ 97 98 100 -1 ]
  //: joint g100 (W) @(2353, 314) /w:[ 29 30 32 -1 ]
  //: joint g74 (Reloj) @(2734, 284) /w:[ 13 14 16 -1 ]
  //: joint g56 (Reloj) @(1008, 284) /w:[ 85 86 88 -1 ]
  FlipFlopD g14 (.Reloj(Reloj), .D(w51), .W(W), .nQ(w53), .Q(w54));   //: @(932, 197) /sz:(40, 40) /sn:0 /p:[ Li0>91 Li1>0 Bi0>91 Ro0<0 Ro1<1 ]
  FlipFlopD g5 (.Reloj(Reloj), .D(w10), .W(W), .nQ(w14), .Q(w13));   //: @(305, 199) /sz:(40, 40) /sn:0 /p:[ Li0>115 Li1>0 Bi0>115 Ro0<0 Ro1<1 ]
  //: joint g95 (W) @(1916, 314) /w:[ 49 50 52 -1 ]
  //: joint g94 (W) @(1825, 314) /w:[ 53 54 56 -1 ]
  //: joint g80 (W) @(428, 314) /w:[ 109 110 112 -1 ]
  //: joint g79 (W) @(338, 314) /w:[ 113 114 116 -1 ]
  //: joint g47 (Reloj) @(116, 284) /w:[ 121 122 124 -1 ]
  assign {w195, w186, w177, w162} = Din; //: CONCAT g44  @(70,41) /sn:0 /R:2 /w:[ 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: joint g105 (W) @(2865, 314) /w:[ 9 10 12 -1 ]
  //: joint g92 (W) @(1574, 314) /w:[ 61 62 64 -1 ]
  //: joint g85 (W) @(962, 314) /w:[ 89 90 92 -1 ]
  //: joint g84 (W) @(772, 314) /w:[ 93 94 96 -1 ]
  assign {w131, w121, w156, w146, w151, w126, w136, w141} = w162; //: CONCAT g36  @(2832,91) /sn:0 /R:1 /w:[ 1 1 1 1 1 1 1 0 1 ] /dr:0 /tp:0 /drp:0
  FlipFlopD g24 (.Reloj(Reloj), .D(w101), .W(W), .nQ(w103), .Q(w104));   //: @(2320, 193) /sz:(40, 40) /sn:0 /p:[ Li0>31 Li1>1 Bi0>31 Ro0<0 Ro1<0 ]
  FlipFlopD g21 (.Reloj(Reloj), .D(w86), .W(W), .nQ(w88), .Q(w89));   //: @(2146, 195) /sz:(40, 40) /sn:0 /p:[ Li0>39 Li1>1 Bi0>39 Ro0<0 Ro1<0 ]
  assign w213 = {w94, w84, w119, w109, w114, w89, w99, w104}; //: CONCAT g41  @(2109,381) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 1 1 1 ] /dr:1 /tp:0 /drp:1
  FlipFlopD g23 (.Reloj(Reloj), .D(w96), .W(W), .nQ(w98), .Q(w99));   //: @(2231, 194) /sz:(40, 40) /sn:0 /p:[ Li0>35 Li1>0 Bi0>35 Ro0<0 Ro1<0 ]
  //: joint g101 (W) @(2517, 314) /w:[ 25 26 28 -1 ]
  //: joint g93 (W) @(1735, 314) /w:[ 57 58 60 -1 ]
  //: joint g81 (W) @(515, 314) /w:[ 105 106 108 -1 ]
  //: joint g60 (Reloj) @(1352, 284) /w:[ 69 70 72 -1 ]
  //: joint g54 (Reloj) @(731, 284) /w:[ 93 94 96 -1 ]
  assign w204 = {w134, w124, w159, w149, w154, w129, w197, w144}; //: CONCAT g40  @(2857,380) /sn:0 /R:3 /w:[ 1 1 1 0 1 0 1 0 1 ] /dr:1 /tp:0 /drp:1
  //: joint g90 (W) @(1402, 314) /w:[ 69 70 72 -1 ]
  //: joint g70 (Reloj) @(2305, 284) /w:[ 29 30 32 -1 ]
  //: joint g46 (Reloj) @(2992, 284) /w:[ 6 8 5 -1 ]
  assign Dout = {w231, w222, w213, w204}; //: CONCAT g45  @(3198,423) /sn:0 /w:[ 0 0 0 0 0 ] /dr:0 /tp:0 /drp:1
  FlipFlopD g35 (.Reloj(Reloj), .D(w156), .W(W), .nQ(w158), .Q(w159));   //: @(2659, 193) /sz:(40, 40) /sn:0 /p:[ Li0>19 Li1>0 Bi0>19 Ro0<0 Ro1<1 ]
  FlipFlopD g26 (.Reloj(Reloj), .D(w111), .W(W), .nQ(w113), .Q(w114));   //: @(2058, 193) /sz:(40, 40) /sn:0 /p:[ Li0>43 Li1>0 Bi0>43 Ro0<0 Ro1<1 ]
  FlipFlopD g22 (.Reloj(Reloj), .D(w91), .W(W), .nQ(w93), .Q(w94));   //: @(1710, 194) /sz:(40, 40) /sn:0 /p:[ Li0>59 Li1>0 Bi0>59 Ro0<0 Ro1<1 ]
  //: IN g0 (Din) @(10,40) /sn:0 /w:[ 0 ]
  //: joint g97 (W) @(2088, 314) /w:[ 41 42 44 -1 ]
  //: joint g82 (W) @(605, 314) /w:[ 101 102 104 -1 ]
  //: joint g66 (Reloj) @(1958, 284) /w:[ 45 46 48 -1 ]
  FlipFlopD g18 (.Reloj(Reloj), .D(w71), .W(W), .nQ(w73), .Q(w74));   //: @(1280, 196) /sz:(40, 40) /sn:0 /p:[ Li0>75 Li1>0 Bi0>75 Ro0<0 Ro1<1 ]
  FlipFlopD g12 (.Reloj(Reloj), .D(w41), .W(W), .nQ(w43), .Q(w44));   //: @(1020, 199) /sz:(40, 40) /sn:0 /p:[ Li0>87 Li1>0 Bi0>87 Ro0<0 Ro1<1 ]
  //: joint g91 (W) @(1482, 314) /w:[ 65 66 68 -1 ]
  FlipFlopD g33 (.Reloj(Reloj), .D(w146), .W(W), .nQ(w148), .Q(w149));   //: @(2748, 192) /sz:(40, 40) /sn:0 /p:[ Li0>15 Li1>0 Bi0>15 Ro0<0 Ro1<0 ]
  FlipFlopD g30 (.Reloj(Reloj), .D(w131), .W(W), .nQ(w133), .Q(w134));   //: @(2486, 192) /sz:(40, 40) /sn:0 /p:[ Li0>27 Li1>0 Bi0>27 Ro0<0 Ro1<0 ]
  //: joint g49 (Reloj) @(292, 284) /w:[ 113 114 116 -1 ]

endmodule
//: /netlistEnd

//: /netlistBegin FlipFlopSR
module FlipFlopSR(nQ, R, S, Reloj, Q);
//: interface  /sz:(134, 64) /bd:[ Li0>R(52/64) Li1>Reloj(32/64) Li2>S(14/64) Ro0<nQ(44/64) Ro1<Q(27/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output Q;    //: /sn:0 {0}(453,103)(545,103)(545,100)(560,100){1}
output nQ;    //: /sn:0 {0}(453,123)(550,123)(550,157)(565,157){1}
input R;    //: /sn:0 {0}(58,157)(154,157)(154,130)(179,130){1}
input Reloj;    //: /sn:0 {0}(56,266)(89,266)(89,238)(104,238){1}
input S;    //: /sn:0 {0}(56,92)(131,92)(131,95)(179,95){1}
wire w7;    //: /sn:0 {0}(287,255)(355,255)(355,111)(370,111){1}
wire w4;    //: /sn:0 {0}(262,104)(273,104)(273,94)(370,94){1}
wire w3;    //: /sn:0 {0}(262,124)(331,124)(331,129)(370,129){1}
wire w0;    //: /sn:0 {0}(179,112)(148,112)(148,264){1}
//: {2}(150,266)(160,266)(160,255)(271,255){3}
//: {4}(146,266)(128,266)(128,238)(120,238){5}
//: enddecls

  _GGNBUF #(2) g4 (.I(Reloj), .Z(w0));   //: @(110,238) /sn:0 /w:[ 1 5 ]
  //: OUT g8 (nQ) @(562,157) /sn:0 /w:[ 1 ]
  //: IN g3 (R) @(56,157) /sn:0 /w:[ 0 ]
  //: IN g2 (S) @(54,92) /sn:0 /w:[ 0 ]
  LatchSR g1 (.C(w7), .R(w3), .S(w4), .nQ(nQ), .Q(Q));   //: @(371, 83) /sz:(81, 64) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Ro0<0 Ro1<0 ]
  //: comment g10 @(266,23) /sn:0
  //: /line:"Flancao ascendente"
  //: /end
  //: IN g6 (Reloj) @(54,266) /sn:0 /w:[ 0 ]
  //: OUT g7 (Q) @(557,100) /sn:0 /w:[ 1 ]
  //: joint g9 (w0) @(148, 266) /w:[ 2 1 4 -1 ]
  _GGNBUF #(2) g5 (.I(w0), .Z(w7));   //: @(277,255) /sn:0 /w:[ 3 0 ]
  LatchSR g0 (.C(w0), .R(R), .S(S), .nQ(w3), .Q(w4));   //: @(180, 84) /sz:(81, 64) /sn:0 /p:[ Li0>0 Li1>1 Li2>1 Ro0<0 Ro1<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FlipFlopT
module FlipFlopT(Q, nQ, Reloj, T);
//: interface  /sz:(106, 65) /bd:[ Li0>Reloj(45/65) Li1>T(25/65) Ro0<nQ(37/65) Ro1<Q(17/65) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output Q;    //: /sn:0 {0}(334,147)(365,147)(365,148)(391,148){1}
//: {2}(395,148)(445,148){3}
//: {4}(393,146)(393,93)(179,93)(179,117)(183,117){5}
//: {6}(393,150)(393,215)(306,215)(306,229)(310,229){7}
output nQ;    //: /sn:0 {0}(172,254)(162,254)(162,284)(385,284)(385,234){1}
//: {2}(387,232)(436,232)(436,236)(447,236){3}
//: {4}(383,232)(374,232)(374,231)(368,231){5}
//: {6}(366,229)(366,163)(301,163)(301,149)(313,149){7}
//: {8}(364,231)(346,231)(346,232)(331,232){9}
input T;    //: /sn:0 {0}(41,125)(98,125){1}
//: {2}(102,125)(147,125)(147,122)(183,122){3}
//: {4}(100,127)(100,249)(172,249){5}
input Reloj;    //: /sn:0 {0}(57,174)(141,174)(141,178)(155,178){1}
//: {2}(157,176)(157,127)(183,127){3}
//: {4}(157,180)(157,244)(172,244){5}
wire w6;    //: /sn:0 {0}(193,249)(295,249)(295,234)(310,234){1}
wire w2;    //: /sn:0 {0}(204,122)(298,122)(298,144)(313,144){1}
//: enddecls

  //: OUT g4 (Q) @(442,148) /sn:0 /w:[ 3 ]
  _GGNOR2 #(4) g8 (.I0(Q), .I1(w6), .Z(nQ));   //: @(321,232) /sn:0 /w:[ 7 1 9 ]
  //: comment g13 @(179,46) /sn:0
  //: /line:"Como pone en internet(no funciona)"
  //: /end
  //: OUT g3 (nQ) @(444,236) /sn:0 /w:[ 3 ]
  //: joint g2 (T) @(100, 125) /w:[ 2 -1 1 4 ]
  //: IN g1 (Reloj) @(55,174) /sn:0 /w:[ 0 ]
  //: joint g11 (nQ) @(366, 231) /w:[ 5 6 8 -1 ]
  //: joint g10 (Q) @(393, 148) /w:[ 2 4 1 6 ]
  _GGAND3 #(8) g6 (.I0(Reloj), .I1(T), .I2(nQ), .Z(w6));   //: @(183,249) /sn:0 /w:[ 5 5 0 0 ]
  _GGNOR2 #(4) g7 (.I0(w2), .I1(nQ), .Z(Q));   //: @(324,147) /sn:0 /w:[ 1 7 0 ]
  //: joint g9 (Reloj) @(157, 178) /w:[ -1 2 1 4 ]
  _GGAND3 #(8) g5 (.I0(Q), .I1(T), .I2(Reloj), .Z(w2));   //: @(194,122) /sn:0 /w:[ 5 3 3 0 ]
  //: IN g0 (T) @(39,125) /sn:0 /w:[ 0 ]
  //: joint g12 (nQ) @(385, 232) /w:[ 2 -1 4 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin ALU
module ALU(Sa, Cero, B, A, C, Overflow);
//: interface  /sz:(129, 64) /bd:[ Ti0>C[2:0](61/129) Li0>A[31:0](19/64) Li1>B[31:0](43/64) Ro0<Cero(31/64) Ro1<Overflow(49/64) Ro2<Sa[31:0](13/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [31:0] A;    //: /sn:0 {0}(#:-133,-78)(-114,-78)(-114,-226)(#:71,-226){1}
supply0 w54;    //: /sn:0 {0}(476,-314)(476,-361){1}
//: {2}(478,-363)(509,-363){3}
//: {4}(476,-365)(476,-372)(509,-372){5}
//: {6}(478,-363)(468,-363)(468,-353)(509,-353){7}
output Cero;    //: /sn:0 {0}(1741,915)(1731,915)(1731,916)(1675,916){1}
output Overflow;    //: /sn:0 {0}(383,2652)(383,2708)(413,2708){1}
output [31:0] Sa;    //: /sn:0 {0}(#:1263,925)(1138,925)(1138,1133){1}
//: {2}(1140,1135)(1325,1135){3}
//: {4}(1136,1135)(#:1034,1135){5}
input [2:0] C;    //: /sn:0 {0}(#:537,2331)(537,2253){1}
//: {2}(539,2251)(716,2251)(716,2169){3}
//: {4}(716,2165)(716,2079){5}
//: {6}(716,2075)(716,1998){7}
//: {8}(716,1994)(716,1913){9}
//: {10}(716,1909)(716,1828){11}
//: {12}(716,1824)(716,1748){13}
//: {14}(716,1744)(716,1661){15}
//: {16}(716,1657)(716,1575){17}
//: {18}(716,1571)(716,1489){19}
//: {20}(716,1485)(716,1416){21}
//: {22}(716,1412)(716,1340){23}
//: {24}(716,1336)(716,1238){25}
//: {26}(716,1234)(716,1151){27}
//: {28}(716,1147)(716,1094){29}
//: {30}(716,1090)(716,992){31}
//: {32}(716,988)(716,898){33}
//: {34}(716,894)(716,826){35}
//: {36}(716,822)(716,741){37}
//: {38}(716,737)(716,657){39}
//: {40}(716,653)(716,561){41}
//: {42}(716,557)(716,461){43}
//: {44}(716,457)(716,373){45}
//: {46}(716,369)(716,284){47}
//: {48}(716,280)(716,197){49}
//: {50}(716,193)(716,140)(717,140)(717,106){51}
//: {52}(717,102)(717,6){53}
//: {54}(717,2)(717,-80){55}
//: {56}(717,-84)(717,-172){57}
//: {58}(717,-176)(717,-277){59}
//: {60}(717,-281)(717,-536)(575,-536){61}
//: {62}(573,-538)(573,-543)(541,-543)(#:541,-546){63}
//: {64}(573,-534)(573,-526)(541,-526)(#:541,-515){65}
//: {66}(715,-279)(431,-279)(431,-257){67}
//: {68}(715,-174)(432,-174)(432,-160){69}
//: {70}(715,-82)(433,-82)(433,-63){71}
//: {72}(715,4)(434,4)(#:434,27){73}
//: {74}(715,104)(435,104)(#:435,118){75}
//: {76}(714,195)(436,195)(#:436,211){77}
//: {78}(714,282)(437,282)(#:437,299){79}
//: {80}(714,371)(438,371)(#:438,393){81}
//: {82}(714,459)(439,459)(#:439,481){83}
//: {84}(714,559)(442,559)(#:442,572){85}
//: {86}(714,655)(509,655)(509,645)(452,645)(#:452,661){87}
//: {88}(714,739)(462,739)(#:462,744){89}
//: {90}(714,824)(444,824)(#:444,829){91}
//: {92}(714,896)(440,896)(#:440,913){93}
//: {94}(714,990)(436,990)(#:436,999){95}
//: {96}(714,1092)(521,1092)(521,1070)(444,1070)(#:444,1082){97}
//: {98}(714,1149)(439,1149)(#:439,1170){99}
//: {100}(714,1236)(459,1236)(#:459,1263){101}
//: {102}(714,1338)(515,1338)(515,1329)(471,1329)(#:471,1343){103}
//: {104}(714,1414)(454,1414)(#:454,1424){105}
//: {106}(714,1487)(451,1487)(#:451,1507){107}
//: {108}(714,1573)(444,1573)(#:444,1592){109}
//: {110}(714,1659)(439,1659)(#:439,1673){111}
//: {112}(714,1746)(451,1746)(#:451,1753){113}
//: {114}(714,1826)(444,1826)(#:444,1839){115}
//: {116}(714,1911)(442,1911)(#:442,1920){117}
//: {118}(714,1996)(429,1996)(#:429,2005){119}
//: {120}(714,2077)(454,2077)(#:454,2093){121}
//: {122}(714,2167)(440,2167)(#:440,2172){123}
//: {124}(535,2251)(461,2251)(#:461,2256){125}
input [31:0] B;    //: /sn:0 {0}(#:-653,763)(#:-290,763){1}
supply0 w49;    //: /sn:0 {0}(467,2432)(441,2432){1}
//: {2}(439,2430)(439,2423)(467,2423){3}
//: {4}(439,2434)(439,2446)(449,2446){5}
//: {6}(451,2444)(451,2442)(467,2442){7}
//: {8}(451,2448)(451,2461){9}
//: {10}(453,2463)(467,2463){11}
//: {12}(451,2465)(451,2498){13}
wire w32;    //: /sn:0 {0}(332,2481)(297,2481){1}
//: {2}(293,2481)(98,2481)(98,2409){3}
//: {4}(100,2407)(110,2407)(110,2412)(292,2412){5}
//: {6}(98,2405)(98,2394){7}
//: {8}(100,2392)(110,2392)(110,2395)(292,2395){9}
//: {10}(98,2390)(98,-71)(77,-71){11}
//: {12}(295,2483)(295,2563)(371,2563)(371,2607){13}
wire w45;    //: /sn:0 {0}(-284,728)(355,728)(355,781)(395,781){1}
wire w73;    //: /sn:0 {0}(1028,1050)(981,1050)(981,331)(459,331){1}
wire w96;    //: /sn:0 {0}(1028,1280)(857,1280)(857,2288)(483,2288){1}
wire w214;    //: /sn:0 {0}(384,1544)(304,1544)(304,818)(-284,818){1}
wire w244;    //: /sn:0 {0}(394,2293)(257,2293)(257,908)(-284,908){1}
wire w122;    //: /sn:0 {0}(398,-98)(398,-79)(370,-79)(370,-70)(398,-70)(398,-63){1}
wire w134;    //: /sn:0 {0}(369,248)(275,248)(275,668)(-284,668){1}
wire w166;    //: /sn:0 {0}(377,866)(350,866)(350,738)(-284,738){1}
wire w203;    //: /sn:0 {0}(419,1424)(419,1415)(437,1415)(437,1405){1}
wire w220;    //: /sn:0 {0}(375,1957)(279,1957)(279,868)(-284,868){1}
wire w141;    //: /sn:0 {0}(403,361)(403,378)(394,378)(394,385)(403,385)(403,393){1}
wire w14;    //: /sn:0 {0}(77,-251)(167,-251)(167,851)(377,851){1}
wire w16;    //: /sn:0 {0}(77,-231)(158,-231)(158,1021)(369,1021){1}
wire w56;    //: /sn:0 {0}(372,1710)(294,1710)(294,838)(-284,838){1}
wire w179;    //: /sn:0 {0}(409,1082)(409,1076)(402,1076)(402,1061){1}
wire w4;    //: /sn:0 {0}(77,-351)(214,-351)(214,-41)(366,-41){1}
wire w19;    //: /sn:0 {0}(392,1285)(144,1285)(144,-201)(77,-201){1}
wire w81;    //: /sn:0 {0}(1028,1130)(943,1130)(943,1031)(458,1031){1}
wire w89;    //: /sn:0 {0}(461,1705)(789,1705)(789,1210)(1028,1210){1}
wire w195;    //: /sn:0 {0}(473,1785)(798,1785)(798,1220)(1028,1220){1}
wire w38;    //: /sn:0 {0}(368,155)(265,155)(265,658)(-284,658){1}
wire w152;    //: /sn:0 {0}(371,430)(301,430)(301,688)(-284,688){1}
wire w3;    //: /sn:0 {0}(77,-361)(218,-361)(218,-138)(365,-138){1}
wire w0;    //: /sn:0 {0}(362,-334)(325,-334)(325,-362){1}
//: {2}(327,-364)(347,-364){3}
//: {4}(325,-366)(325,-379){5}
//: {6}(327,-381)(347,-381){7}
//: {8}(323,-381)(77,-381){9}
wire w151;    //: /sn:0 {0}(377,1629)(298,1629)(298,828)(-284,828){1}
wire w128;    //: /sn:0 {0}(1269,1060)(1609,1060)(1609,984)(1654,984){1}
wire w127;    //: /sn:0 {0}(1269,1050)(1599,1050)(1599,979)(1654,979){1}
wire w120;    //: /sn:0 {0}(1028,1000)(1000,1000)(1000,-128)(454,-128){1}
wire w233;    //: /sn:0 {0}(405,2172)(405,2165)(420,2165)(420,2155){1}
wire w240;    //: /sn:0 {0}(1028,1270)(846,1270)(846,2204)(462,2204){1}
wire w133;    //: /sn:0 {0}(-284,708)(320,708)(320,609)(375,609){1}
wire w104;    //: /sn:0 {0}(396,-288)(396,-274)(385,-274)(385,-266)(396,-266)(396,-257){1}
wire w111;    //: /sn:0 {0}(368,-378)(428,-378)(428,-403)(509,-403){1}
wire w168;    //: /sn:0 {0}(1028,1110)(954,1110)(954,861)(466,861){1}
wire w204;    //: /sn:0 {0}(1028,1170)(750,1170)(750,1375)(493,1375){1}
wire w75;    //: /sn:0 {0}(1028,1070)(973,1070)(973,513)(461,513){1}
wire w209;    //: /sn:0 {0}(416,1507)(416,1495)(420,1495)(420,1486){1}
wire w67;    //: /sn:0 {0}(1028,990)(1005,990)(1005,-225)(453,-225){1}
wire w119;    //: /sn:0 {0}(400,118)(400,106)(387,106)(387,97)(400,97)(400,89){1}
wire w90;    //: /sn:0 {0}(1269,910)(1513,910)(1513,909)(1654,909){1}
wire w215;    //: /sn:0 {0}(409,1592)(409,1574)(417,1574)(417,1569){1}
wire w156;    //: /sn:0 {0}(1028,1090)(965,1090)(965,693)(474,693){1}
wire w167;    //: /sn:0 {0}(405,913)(405,904)(396,904)(396,896)(410,896)(410,891){1}
wire w41;    //: /sn:0 {0}(313,2415)(387,2415)(387,2404)(467,2404){1}
wire w36;    //: /sn:0 {0}(366,-26)(252,-26)(252,638)(-284,638){1}
wire w20;    //: /sn:0 {0}(77,-191)(139,-191)(139,1365)(404,1365){1}
wire w23;    //: /sn:0 {0}(377,1614)(129,1614)(129,-161)(77,-161){1}
wire w124;    //: /sn:0 {0}(1028,1020)(992,1020)(992,59)(456,59){1}
wire w174;    //: /sn:0 {0}(1028,1120)(949,1120)(949,945)(462,945){1}
wire w82;    //: /sn:0 {0}(1028,1140)(939,1140)(939,1114)(466,1114){1}
wire w126;    //: /sn:0 {0}(1028,1010)(996,1010)(996,-31)(455,-31){1}
wire w74;    //: /sn:0 {0}(1028,1060)(977,1060)(977,425)(460,425){1}
wire w125;    //: /sn:0 {0}(399,-1)(399,13)(371,13)(371,19)(399,19)(399,27){1}
wire w91;    //: /sn:0 {0}(466,1871)(806,1871)(806,1230)(1028,1230){1}
wire w35;    //: /sn:0 {0}(365,-123)(247,-123)(247,628)(-284,628){1}
wire w8;    //: /sn:0 {0}(77,-311)(195,-311)(195,321)(370,321){1}
wire w103;    //: /sn:0 {0}(551,-509)(551,-467)(552,-467)(552,-411){1}
wire w101;    //: /sn:0 {0}(1269,970)(1542,970)(1542,939)(1654,939){1}
wire w192;    //: /sn:0 {0}(461,1202)(724,1202)(724,1150)(1028,1150){1}
wire w71;    //: /sn:0 {0}(1028,1030)(988,1030)(988,150)(457,150){1}
wire w202;    //: /sn:0 {0}(404,1380)(313,1380)(313,798)(-284,798){1}
wire w238;    //: /sn:0 {0}(373,2209)(261,2209)(261,898)(-284,898){1}
wire w22;    //: /sn:0 {0}(384,1529)(133,1529)(133,-171)(77,-171){1}
wire w17;    //: /sn:0 {0}(377,1104)(153,1104)(153,-221)(77,-221){1}
wire w117;    //: /sn:0 {0}(1269,1010)(1563,1010)(1563,959)(1654,959){1}
wire w53;    //: /sn:0 {0}(387,1461)(308,1461)(308,808)(-284,808){1}
wire w84;    //: /sn:0 {0}(1028,1160)(739,1160)(739,1295)(481,1295){1}
wire w172;    //: /sn:0 {0}(-284,748)(344,748)(344,950)(373,950){1}
wire w211;    //: /sn:0 {0}(407,1920)(407,1908)(410,1908)(410,1901){1}
wire w228;    //: /sn:0 {0}(1028,1250)(823,1250)(823,2037)(451,2037){1}
wire w12;    //: /sn:0 {0}(385,683)(177,683)(177,-271)(77,-271){1}
wire w113;    //: /sn:0 {0}(397,-195)(397,-180)(383,-180)(383,-172)(397,-172)(397,-160){1}
wire w44;    //: /sn:0 {0}(-284,718)(326,718)(326,698)(385,698){1}
wire w2;    //: /sn:0 {0}(396,-350)(396,-462){1}
//: {2}(398,-464)(528,-464){3}
//: {4}(530,-466)(530,-496)(531,-496)(531,-509){5}
//: {6}(530,-462)(530,-411){7}
//: {8}(394,-464)(284,-464)(284,-353)(309,-353)(309,-330){9}
wire w115;    //: /sn:0 {0}(1269,990)(1554,990)(1554,949)(1654,949){1}
wire w83;    //: /sn:0 {0}(1269,870)(1548,870)(1548,889)(1654,889){1}
wire w77;    //: /sn:0 {0}(1269,850)(1569,850)(1569,879)(1654,879){1}
wire w226;    //: /sn:0 {0}(362,2042)(273,2042)(273,878)(-284,878){1}
wire w78;    //: /sn:0 {0}(1028,1100)(960,1100)(960,776)(484,776){1}
wire w10;    //: /sn:0 {0}(372,503)(186,503)(186,-291)(77,-291){1}
wire w27;    //: /sn:0 {0}(375,1942)(114,1942)(114,-121)(77,-121){1}
wire w190;    //: /sn:0 {0}(372,1207)(326,1207)(326,778)(-284,778){1}
wire w95;    //: /sn:0 {0}(1269,940)(1528,940)(1528,924)(1654,924){1}
wire w52;    //: /sn:0 {0}(1028,1290)(869,1290)(869,2426)(521,2426){1}
wire w86;    //: /sn:0 {0}(1028,1180)(762,1180)(762,1456)(476,1456){1}
wire w80;    //: /sn:0 {0}(213,2538)(142,2538){1}
//: {2}(138,2538)(97,2538){3}
//: {4}(93,2538)(-18,2538)(-18,2412){5}
//: {6}(-16,2410)(-6,2410)(-6,2417)(292,2417){7}
//: {8}(-18,2408)(-18,918)(-284,918){9}
//: {10}(-20,2410)(-30,2410)(-30,2400)(292,2400){11}
//: {12}(95,2540)(95,2588)(392,2588)(392,2607){13}
//: {14}(140,2540)(140,2556)(157,2556){15}
wire w29;    //: /sn:0 {0}(387,2115)(107,2115)(107,-101)(77,-101){1}
wire w155;    //: /sn:0 {0}(427,744)(427,735)(418,735)(418,723){1}
wire w178;    //: /sn:0 {0}(369,1036)(338,1036)(338,758)(-284,758){1}
wire w50;    //: /sn:0 {0}(1269,780)(1628,780)(1628,844)(1654,844){1}
wire w147;    //: /sn:0 {0}(407,572)(407,562)(399,562)(399,553)(405,553)(405,543){1}
wire w42;    //: /sn:0 {0}(-284,698)(311,698)(311,518)(372,518){1}
wire w6;    //: /sn:0 {0}(77,-331)(204,-331)(204,140)(368,140){1}
wire w93;    //: /sn:0 {0}(1654,914)(1517,914)(1517,920)(1269,920){1}
wire w7;    //: /sn:0 {0}(77,-321)(199,-321)(199,233)(369,233){1}
wire w99;    //: /sn:0 {0}(1269,960)(1536,960)(1536,934)(1654,934){1}
wire w175;    //: /sn:0 {0}(416,1753)(416,1744)(405,1744)(405,1735){1}
wire w112;    //: /sn:0 {0}(77,-371)(221,-371)(221,-235)(364,-235){1}
wire w61;    //: /sn:0 {0}(387,2130)(267,2130)(267,888)(-284,888){1}
wire w135;    //: /sn:0 {0}(402,299)(402,286)(394,286)(394,279)(402,279)(402,273){1}
wire w15;    //: /sn:0 {0}(373,935)(163,935)(163,-241)(77,-241){1}
wire w216;    //: /sn:0 {0}(473,1539)(771,1539)(771,1190)(1028,1190){1}
wire w69;    //: /sn:0 {0}(1269,820)(1591,820)(1591,864)(1654,864){1}
wire w239;    //: /sn:0 {0}(426,2256)(426,2244)(406,2244)(406,2234){1}
wire w207;    //: /sn:0 {0}(377,1876)(283,1876)(283,858)(-284,858){1}
wire w51;    //: /sn:0 {0}(392,1300)(319,1300)(319,788)(-284,788){1}
wire w109;    //: /sn:0 {0}(364,-220)(242,-220)(242,618)(-284,618){1}
wire w129;    //: /sn:0 {0}(401,211)(401,193)(391,193)(391,185)(401,185)(401,180){1}
wire w114;    //: /sn:0 {0}(1269,980)(1548,980)(1548,944)(1654,944){1}
wire w97;    //: /sn:0 {0}(1269,950)(1532,950)(1532,929)(1654,929){1}
wire w64;    //: /sn:0 {0}(1269,810)(1599,810)(1599,859)(1654,859){1}
wire w66;    //: /sn:0 {0}(563,-369)(1010,-369)(1010,980)(1028,980){1}
wire w37;    //: /sn:0 {0}(367,64)(257,64)(257,648)(-284,648){1}
wire w245;    //: /sn:0 {0}(427,2318)(427,2374)(366,2374)(366,2465){1}
wire w63;    //: /sn:0 {0}(1269,800)(1608,800)(1608,854)(1654,854){1}
wire w34;    //: /sn:0 {0}(537,2337)(537,2365)(499,2365)(499,2384){1}
wire w234;    //: /sn:0 {0}(1028,1260)(834,1260)(834,2125)(476,2125){1}
wire w159;    //: /sn:0 {0}(466,1624)(780,1624)(780,1200)(1028,1200){1}
wire w21;    //: /sn:0 {0}(77,-181)(136,-181)(136,1446)(387,1446){1}
wire w76;    //: /sn:0 {0}(1028,1080)(969,1080)(969,604)(464,604){1}
wire w102;    //: /sn:0 {0}(541,-509)(541,-411){1}
wire w157;    //: /sn:0 {0}(404,1673)(404,1662)(410,1662)(410,1654){1}
wire w43;    //: /sn:0 {0}(1269,770)(1639,770)(1639,839)(1654,839){1}
wire w87;    //: /sn:0 {0}(1269,890)(1532,890)(1532,899)(1654,899){1}
wire w31;    //: /sn:0 {0}(394,2278)(101,2278)(101,-81)(77,-81){1}
wire w100;    //: /sn:0 {0}(431,-321)(455,-321)(455,-340){1}
//: {2}(457,-342)(509,-342){3}
//: {4}(455,-344)(455,-383)(509,-383){5}
wire w28;    //: /sn:0 {0}(362,2027)(111,2027)(111,-111)(77,-111){1}
wire w130;    //: /sn:0 {0}(1269,1070)(1625,1070)(1625,989)(1654,989){1}
wire w24;    //: /sn:0 {0}(77,-151)(126,-151)(126,1695)(372,1695){1}
wire w184;    //: /sn:0 {0}(377,1119)(332,1119)(332,768)(-284,768){1}
wire w161;    //: /sn:0 {0}(409,829)(409,815)(428,815)(428,806){1}
wire w1;    //: /sn:0 {0}(547,2337)(547,2371)(510,2371)(510,2384){1}
wire w140;    //: /sn:0 {0}(370,336)(289,336)(289,678)(-284,678){1}
wire w221;    //: /sn:0 {0}(394,2005)(394,1989)(408,1989)(408,1982){1}
wire w25;    //: /sn:0 {0}(77,-141)(123,-141)(123,1775)(384,1775){1}
wire w98;    //: /sn:0 {0}(288,-301)(256,-301){1}
wire w65;    //: /sn:0 {0}(467,2453)(448,2453){1}
//: {2}(444,2453)(426,2453){3}
//: {4}(424,2451)(424,2412)(467,2412){5}
//: {6}(424,2455)(424,2492){7}
//: {8}(422,2494)(401,2494){9}
//: {10}(424,2496)(424,2558)(414,2558)(414,2607){11}
//: {12}(446,2455)(446,2488)(437,2488)(437,2526)(620,2526)(620,-317)(499,-317)(499,-332)(509,-332){13}
wire w227;    //: /sn:0 {0}(419,2093)(419,2079)(395,2079)(395,2067){1}
wire w116;    //: /sn:0 {0}(1269,1000)(1559,1000)(1559,954)(1654,954){1}
wire w18;    //: /sn:0 {0}(372,1192)(148,1192)(148,-211)(77,-211){1}
wire w92;    //: /sn:0 {0}(1028,1240)(815,1240)(815,1952)(464,1952){1}
wire w40;    //: /sn:0 {0}(313,2398)(445,2398)(445,2392)(467,2392){1}
wire w118;    //: /sn:0 {0}(1269,1020)(1568,1020)(1568,964)(1654,964){1}
wire w121;    //: /sn:0 {0}(1269,1030)(1575,1030)(1575,969)(1654,969){1}
wire w30;    //: /sn:0 {0}(373,2194)(104,2194)(104,-91)(77,-91){1}
wire w68;    //: /sn:0 {0}(173,2556)(213,2556){1}
wire w59;    //: /sn:0 {0}(366,2527)(366,2542){1}
wire w123;    //: /sn:0 {0}(1269,1040)(1586,1040)(1586,974)(1654,974){1}
wire w185;    //: /sn:0 {0}(404,1170)(404,1155)(410,1155)(410,1144){1}
wire w62;    //: /sn:0 {0}(1269,790)(1616,790)(1616,849)(1654,849){1}
wire w85;    //: /sn:0 {0}(1269,880)(1540,880)(1540,894)(1654,894){1}
wire w173;    //: /sn:0 {0}(401,999)(401,986)(406,986)(406,975){1}
wire w136;    //: /sn:0 {0}(1028,1040)(985,1040)(985,243)(458,243){1}
wire w57;    //: /sn:0 {0}(384,1790)(288,1790)(288,848)(-284,848){1}
wire w11;    //: /sn:0 {0}(375,594)(182,594)(182,-281)(77,-281){1}
wire w137;    //: /sn:0 {0}(417,661)(417,650)(408,650)(408,634){1}
wire w197;    //: /sn:0 {0}(436,1343)(436,1335)(425,1335)(425,1325){1}
wire w105;    //: /sn:0 {0}(330,-312)(362,-312){1}
wire w110;    //: /sn:0 {0}(368,-361)(440,-361)(440,-391)(509,-391){1}
wire w193;    //: /sn:0 {0}(409,1839)(409,1826)(417,1826)(417,1815){1}
wire w70;    //: /sn:0 {0}(1269,830)(1584,830)(1584,869)(1654,869){1}
wire w13;    //: /sn:0 {0}(395,766)(172,766)(172,-261)(77,-261){1}
wire w72;    //: /sn:0 {0}(1269,840)(1577,840)(1577,874)(1654,874){1}
wire w88;    //: /sn:0 {0}(1269,900)(1523,900)(1523,904)(1654,904){1}
wire w94;    //: /sn:0 {0}(1654,919)(1524,919)(1524,930)(1269,930){1}
wire w191;    //: /sn:0 {0}(424,1263)(424,1243)(405,1243)(405,1232){1}
wire w33;    //: /sn:0 {0}(347,-376)(307,-376){1}
//: {2}(303,-376)(129,-376)(129,-326){3}
//: {4}(131,-324)(226,-324){5}
//: {6}(230,-324)(259,-324)(259,-319)(288,-319){7}
//: {8}(228,-322)(228,-301)(240,-301){9}
//: {10}(127,-324)(97,-324)(97,-426)(-260,-426)(-260,608)(-284,608){11}
//: {12}(305,-374)(305,-359)(347,-359){13}
wire w5;    //: /sn:0 {0}(77,-341)(209,-341)(209,49)(367,49){1}
wire w143;    //: /sn:0 {0}(404,481)(404,470)(393,470)(393,464)(404,464)(404,455){1}
wire w131;    //: /sn:0 {0}(1269,1080)(1639,1080)(1639,994)(1654,994){1}
wire w9;    //: /sn:0 {0}(77,-301)(191,-301)(191,415)(371,415){1}
wire w79;    //: /sn:0 {0}(1269,860)(1560,860)(1560,884)(1654,884){1}
wire w26;    //: /sn:0 {0}(377,1861)(118,1861)(118,-131)(77,-131){1}
wire w39;    //: /sn:0 {0}(234,2527)(234,2452)(276,2452){1}
//: {2}(280,2452)(341,2452)(341,2359)(486,2359){3}
//: {4}(490,2359)(527,2359)(527,2337){5}
//: {6}(488,2361)(488,2384){7}
//: {8}(278,2454)(278,2571)(349,2571)(349,2607){9}
wire w55;    //: /sn:0 {0}(255,2545)(317,2545)(317,2503)(332,2503){1}
//: enddecls

  //: OUT g4 (Sa) @(1322,1135) /sn:0 /w:[ 3 ]
  ALU1bit g8 (.AcarreoE(w104), .C(C), .A(w112), .B(w109), .AcarreoS(w113), .Sa(w67));   //: @(365, -256) /sz:(87, 60) /sn:0 /p:[ Ti0>1 Ti1>67 Li0>1 Li1>0 Bo0<0 Ro0<1 ]
  //: GROUND g140 (w54) @(476,-308) /sn:0 /w:[ 0 ]
  //: comment g58 @(360,1750) /sn:0
  //: /line:"24"
  //: /end
  //: comment g55 @(333,2005) /sn:0
  //: /line:"27"
  //: /end
  ALU1bit g37 (.C(C), .AcarreoE(w179), .B(w184), .A(w17), .AcarreoS(w185), .Sa(w82));   //: @(378, 1083) /sz:(87, 60) /sn:0 /p:[ Ti0>97 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<1 ]
  //: joint g13 (w0) @(325, -364) /w:[ 2 4 -1 1 ]
  //: OUT g139 (Cero) @(1738,915) /sn:0 /w:[ 0 ]
  //: joint g112 (w80) @(95, 2538) /w:[ 3 -1 4 12 ]
  //: joint g76 (C) @(716, 990) /w:[ -1 32 94 31 ]
  //: joint g111 (w32) @(295, 2481) /w:[ 1 -1 2 12 ]
  //: IN g1 (B) @(-655,763) /sn:0 /w:[ 0 ]
  //: joint g64 (C) @(717, -82) /w:[ -1 56 70 55 ]
  //: joint g11 (w0) @(325, -381) /w:[ 6 -1 8 5 ]
  //: comment g130 @(363,1155) /sn:0
  //: /line:"17"
  //: /end
  //: comment g121 @(362,385) /sn:0
  //: /line:"8"
  //: /end
  ALU1bit g50 (.C(C), .AcarreoE(w233), .B(w238), .A(w30), .AcarreoS(w239), .Sa(w240));   //: @(374, 2173) /sz:(87, 60) /sn:0 /p:[ Ti0>123 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<1 ]
  ALU1bit g28 (.C(C), .AcarreoE(w135), .B(w140), .A(w8), .AcarreoS(w141), .Sa(w73));   //: @(371, 300) /sz:(87, 60) /sn:0 /p:[ Ti0>79 Ti1>0 Li0>0 Li1>1 Bo0<0 Ro0<1 ]
  //: comment g132 @(390,1335) /sn:0
  //: /line:"19"
  //: /end
  Mux1 g19 (.C(w2), .E0(w33), .E1(w98), .Sal(w105));   //: @(289, -329) /sz:(40, 40) /sn:0 /p:[ Ti0>9 Li0>7 Li1>0 Ro0<0 ]
  //: comment g113 @(345,-295) /sn:0
  //: /line:"0"
  //: /end
  ALU1bit g38 (.C(C), .AcarreoE(w185), .B(w190), .A(w18), .AcarreoS(w191), .Sa(w192));   //: @(373, 1171) /sz:(87, 60) /sn:0 /p:[ Ti0>99 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<0 ]
  Suma g6 (.AcarreoE(w2), .B(w105), .A(w0), .AcarreoS(w104), .Suma(w100));   //: @(363, -349) /sz:(67, 60) /sn:0 /p:[ Ti0>0 Li0>1 Li1>0 Bo0<0 Ro0<0 ]
  //: comment g115 @(355,-172) /sn:0
  //: /line:"2"
  //: /end
  //: comment g53 @(339,2178) /sn:0
  //: /line:"29"
  //: /end
  Mux3 g7 (.C0(w103), .C1(w102), .C2(w2), .E0(w111), .E1(w110), .E2(w100), .E3(w54), .E4(w54), .E5(w54), .E6(w100), .E7(w65), .Sal(w66));   //: @(510, -410) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>7 Li0>1 Li1>1 Li2>5 Li3>5 Li4>3 Li5>7 Li6>3 Li7>13 Ro0<0 ]
  //: joint g75 (C) @(716, 896) /w:[ -1 34 92 33 ]
  //: comment g135 @(392,2437) /sn:0
  //: /line:"31"
  //: /end
  ALU1bit g31 (.C(C), .AcarreoE(w147), .B(w133), .A(w11), .AcarreoS(w137), .Sa(w76));   //: @(376, 573) /sz:(87, 60) /sn:0 /p:[ Ti0>85 Ti1>0 Li0>1 Li1>0 Bo0<1 Ro0<1 ]
  //: joint g20 (w2) @(396, -464) /w:[ 2 -1 8 1 ]
  //: comment g124 @(375,658) /sn:0
  //: /line:"11"
  //: /end
  ALU1bit g39 (.C(C), .AcarreoE(w191), .B(w51), .A(w19), .AcarreoS(w197), .Sa(w84));   //: @(393, 1264) /sz:(87, 60) /sn:0 /p:[ Ti0>101 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<1 ]
  //: joint g68 (C) @(716, 282) /w:[ -1 48 78 47 ]
  ALU1bit g48 (.C(C), .AcarreoE(w221), .B(w226), .A(w28), .AcarreoS(w227), .Sa(w228));   //: @(363, 2006) /sz:(87, 60) /sn:0 /p:[ Ti0>119 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<1 ]
  ALU1bit g29 (.C(C), .AcarreoE(w143), .B(w42), .A(w10), .AcarreoS(w147), .Sa(w75));   //: @(373, 482) /sz:(87, 60) /sn:0 /p:[ Ti0>83 Ti1>0 Li0>1 Li1>0 Bo0<1 Ro0<1 ]
  ALU1bit g25 (.C(C), .AcarreoE(w125), .B(w37), .A(w5), .AcarreoS(w119), .Sa(w124));   //: @(368, 28) /sz:(87, 60) /sn:0 /p:[ Ti0>73 Ti1>1 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  assign {w2, w102, w103} = C; //: CONCAT g17  @(541,-514) /sn:0 /R:1 /w:[ 5 0 0 65 ] /dr:0 /tp:0 /drp:0
  //: joint g106 (w80) @(-18, 2410) /w:[ 6 8 10 5 ]
  //: comment g52 @(370,2262) /sn:0
  //: /line:"30"
  //: /end
  Overflow g107 (.A31(w32), .B31(w80), .R(w39), .SiSa(w65), .Sa(Overflow));   //: @(329, 2608) /sz:(111, 43) /sn:0 /p:[ Ti0>13 Ti1>13 Ti2>9 Ti3>11 Bo0<0 ]
  //: joint g83 (C) @(716, 1573) /w:[ -1 18 108 17 ]
  //: joint g100 (w39) @(488, 2359) /w:[ 4 -1 3 6 ]
  _GGNBUF #(2) g14 (.I(w33), .Z(w98));   //: @(246,-301) /sn:0 /w:[ 9 1 ]
  ALU1bit g47 (.C(C), .AcarreoE(w211), .B(w220), .A(w27), .AcarreoS(w221), .Sa(w92));   //: @(376, 1921) /sz:(87, 60) /sn:0 /p:[ Ti0>117 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<1 ]
  ALU1bit g44 (.C(C), .AcarreoE(w157), .B(w56), .A(w24), .AcarreoS(w175), .Sa(w89));   //: @(373, 1674) /sz:(87, 60) /sn:0 /p:[ Ti0>111 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<0 ]
  //: joint g80 (C) @(716, 1338) /w:[ -1 24 102 23 ]
  _GGAND2 #(6) g94 (.I0(w32), .I1(w80), .Z(w40));   //: @(303,2398) /sn:0 /w:[ 9 11 0 ]
  //: joint g105 (w80) @(140, 2538) /w:[ 1 -1 2 14 ]
  //: joint g21 (w33) @(129, -324) /w:[ 4 3 10 -1 ]
  //: joint g84 (C) @(716, 1659) /w:[ -1 16 110 15 ]
  //: joint g141 (w54) @(476, -363) /w:[ 2 4 6 1 ]
  ALU1bit g41 (.C(C), .AcarreoE(w203), .B(w53), .A(w21), .AcarreoS(w209), .Sa(w86));   //: @(388, 1425) /sz:(87, 60) /sn:0 /p:[ Ti0>105 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  ALU1bit g23 (.AcarreoE(w113), .C(C), .A(w3), .B(w35), .AcarreoS(w122), .Sa(w120));   //: @(366, -159) /sz:(87, 60) /sn:0 /p:[ Ti0>1 Ti1>69 Li0>1 Li1>0 Bo0<0 Ro0<1 ]
  //: comment g54 @(344,2094) /sn:0
  //: /line:"28"
  //: /end
  ALU1bit g40 (.C(C), .AcarreoE(w197), .B(w202), .A(w20), .AcarreoS(w203), .Sa(w204));   //: @(405, 1344) /sz:(87, 60) /sn:0 /p:[ Ti0>103 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  Mux1 g93 (.C(w39), .E1(w68), .E0(w80), .Sal(w55));   //: @(214, 2528) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Li0>1 Li1>0 Ro0<0 ]
  //: comment g116 @(356,-74) /sn:0
  //: /line:"3"
  //: /end
  //: comment g123 @(363,565) /sn:0
  //: /line:"10"
  //: /end
  ALU1bit g46 (.C(C), .AcarreoE(w193), .B(w207), .A(w26), .AcarreoS(w211), .Sa(w91));   //: @(378, 1840) /sz:(87, 60) /sn:0 /p:[ Ti0>115 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<0 ]
  ALU1bit g26 (.C(C), .AcarreoE(w119), .B(w38), .A(w6), .AcarreoS(w129), .Sa(w71));   //: @(369, 119) /sz:(87, 60) /sn:0 /p:[ Ti0>75 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  //: IN g0 (A) @(-135,-78) /sn:0 /w:[ 0 ]
  //: joint g90 (C) @(716, 2167) /w:[ -1 4 122 3 ]
  //: joint g82 (C) @(716, 1487) /w:[ -1 20 106 19 ]
  assign {w131, w130, w128, w127, w123, w121, w118, w117, w116, w115, w114, w101, w99, w97, w95, w94, w93, w90, w88, w87, w85, w83, w79, w77, w72, w70, w69, w64, w63, w62, w50, w43} = Sa; //: CONCAT g136  @(1264,925) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /dr:0 /tp:0 /drp:0
  //: comment g128 @(364,983) /sn:0
  //: /line:"15"
  //: /end
  ALU1bit g33 (.C(C), .AcarreoE(w155), .B(w45), .A(w13), .AcarreoS(w161), .Sa(w78));   //: @(396, 745) /sz:(87, 60) /sn:0 /p:[ Ti0>89 Ti1>0 Li0>1 Li1>0 Bo0<1 Ro0<1 ]
  Mux3 g91 (.C2(w39), .C1(w34), .C0(w1), .E7(w49), .E6(w65), .E5(w49), .E4(w49), .E3(w49), .E2(w65), .E1(w41), .E0(w40), .Sal(w52));   //: @(468, 2385) /sz:(52, 85) /sn:0 /p:[ Ti0>7 Ti1>1 Ti2>1 Li0>11 Li1>0 Li2>7 Li3>0 Li4>3 Li5>5 Li6>1 Li7>1 Ro0<1 ]
  ALU1bit g49 (.C(C), .AcarreoE(w227), .B(w61), .A(w29), .AcarreoS(w233), .Sa(w234));   //: @(388, 2094) /sz:(87, 60) /sn:0 /p:[ Ti0>121 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<1 ]
  _GGNOR32 #(64) g137 (.I0(w43), .I1(w50), .I2(w62), .I3(w63), .I4(w64), .I5(w69), .I6(w70), .I7(w72), .I8(w77), .I9(w79), .I10(w83), .I11(w85), .I12(w87), .I13(w88), .I14(w90), .I15(w93), .I16(w94), .I17(w95), .I18(w97), .I19(w99), .I20(w101), .I21(w114), .I22(w115), .I23(w116), .I24(w117), .I25(w118), .I26(w121), .I27(w123), .I28(w127), .I29(w128), .I30(w130), .I31(w131), .Z(Cero));   //: @(1665,916) /sn:0 /w:[ 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ]
  //: joint g61 (C) @(573, -536) /w:[ 61 62 -1 64 ]
  ALU1bit g51 (.C(C), .AcarreoE(w239), .B(w244), .A(w31), .AcarreoS(w245), .Sa(w96));   //: @(395, 2257) /sz:(87, 60) /sn:0 /p:[ Ti0>125 Ti1>0 Li0>0 Li1>0 Bo0<0 Ro0<1 ]
  ALU1bit g34 (.C(C), .AcarreoE(w161), .B(w166), .A(w14), .AcarreoS(w167), .Sa(w168));   //: @(378, 830) /sz:(87, 60) /sn:0 /p:[ Ti0>91 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  assign {w80, w244, w238, w61, w226, w220, w207, w57, w56, w151, w214, w53, w202, w51, w190, w184, w178, w172, w166, w45, w44, w133, w42, w152, w140, w134, w38, w37, w36, w35, w109, w33} = B; //: CONCAT g3  @(-289,763) /sn:0 /R:2 /w:[ 9 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1 11 1 ] /dr:0 /tp:0 /drp:0
  //: joint g86 (C) @(716, 1826) /w:[ -1 12 114 11 ]
  //: joint g89 (C) @(716, 2077) /w:[ -1 6 120 5 ]
  assign {w32, w31, w30, w29, w28, w27, w26, w25, w24, w23, w22, w21, w20, w19, w18, w17, w16, w15, w14, w13, w12, w11, w10, w9, w8, w7, w6, w5, w4, w3, w112, w0} = A; //: CONCAT g2  @(72,-226) /sn:0 /R:2 /w:[ 11 1 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 9 1 ] /dr:0 /tp:0 /drp:0
  //: joint g65 (C) @(717, 4) /w:[ -1 54 72 53 ]
  //: joint g77 (C) @(716, 1092) /w:[ -1 30 96 29 ]
  //: joint g110 (w65) @(424, 2494) /w:[ -1 7 8 10 ]
  //: comment g59 @(355,1673) /sn:0
  //: /line:"23"
  //: /end
  //: joint g72 (C) @(716, 655) /w:[ -1 40 86 39 ]
  assign {w39, w34, w1} = C; //: CONCAT g98  @(537,2332) /sn:0 /R:1 /w:[ 5 0 0 0 ] /dr:0 /tp:0 /drp:0
  //: joint g99 (C) @(537, 2251) /w:[ 2 -1 124 1 ]
  //: IN g16 (C) @(541,-548) /sn:0 /R:3 /w:[ 63 ]
  //: joint g96 (w65) @(424, 2453) /w:[ 3 4 -1 6 ]
  //: joint g103 (w32) @(98, 2392) /w:[ 8 10 -1 7 ]
  //: comment g122 @(363,473) /sn:0
  //: /line:"9"
  //: /end
  _GGOR2 #(6) g10 (.I0(w0), .I1(w33), .Z(w110));   //: @(358,-361) /sn:0 /w:[ 3 13 0 ]
  //: joint g78 (C) @(716, 1149) /w:[ -1 28 98 27 ]
  //: joint g87 (C) @(716, 1911) /w:[ -1 10 116 9 ]
  //: comment g129 @(364,1074) /sn:0
  //: /line:"16"
  //: /end
  ALU1bit g32 (.C(C), .AcarreoE(w137), .B(w44), .A(w12), .AcarreoS(w155), .Sa(w156));   //: @(386, 662) /sz:(87, 60) /sn:0 /p:[ Ti0>87 Ti1>0 Li0>1 Li1>0 Bo0<1 Ro0<1 ]
  ALU1bit g27 (.C(C), .AcarreoE(w129), .B(w134), .A(w7), .AcarreoS(w135), .Sa(w136));   //: @(370, 212) /sz:(87, 60) /sn:0 /p:[ Ti0>77 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  //: joint g102 (w65) @(446, 2453) /w:[ 1 -1 2 12 ]
  //: joint g143 (w49) @(451, 2446) /w:[ -1 6 5 8 ]
  //: joint g69 (C) @(716, 371) /w:[ -1 46 80 45 ]
  //: comment g57 @(344,1839) /sn:0
  //: /line:"25"
  //: /end
  _GGAND2 #(6) g9 (.I0(w0), .I1(w33), .Z(w111));   //: @(358,-378) /sn:0 /w:[ 7 0 0 ]
  //: comment g119 @(357,206) /sn:0
  //: /line:"6"
  //: /end
  //: joint g142 (w49) @(451, 2463) /w:[ 10 9 -1 12 ]
  //: joint g15 (w100) @(455, -342) /w:[ 2 4 -1 1 ]
  //: joint g71 (C) @(716, 559) /w:[ -1 42 84 41 ]
  //: comment g131 @(379,1252) /sn:0
  //: /line:"18"
  //: /end
  //: joint g67 (C) @(716, 195) /w:[ -1 50 76 49 ]
  //: comment g127 @(365,901) /sn:0
  //: /line:"14"
  //: /end
  ALU1bit g43 (.C(C), .AcarreoE(w215), .B(w151), .A(w23), .AcarreoS(w157), .Sa(w159));   //: @(378, 1593) /sz:(87, 60) /sn:0 /p:[ Ti0>109 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<0 ]
  //: joint g104 (w32) @(98, 2407) /w:[ 4 6 -1 3 ]
  //: joint g62 (C) @(717, -279) /w:[ -1 60 66 59 ]
  //: joint g73 (C) @(716, 739) /w:[ -1 38 88 37 ]
  //: joint g88 (C) @(716, 1996) /w:[ -1 8 118 7 ]
  //: joint g138 (Sa) @(1138, 1135) /w:[ 2 1 4 -1 ]
  ALU1bit g42 (.C(C), .AcarreoE(w209), .B(w214), .A(w22), .AcarreoS(w215), .Sa(w216));   //: @(385, 1508) /sz:(87, 60) /sn:0 /p:[ Ti0>107 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<0 ]
  //: joint g63 (C) @(717, -174) /w:[ -1 58 68 57 ]
  //: joint g74 (C) @(716, 824) /w:[ -1 36 90 35 ]
  //: joint g109 (w39) @(278, 2452) /w:[ 2 -1 1 8 ]
  //: comment g133 @(374,1410) /sn:0
  //: /line:"20"
  //: /end
  //: comment g56 @(346,1923) /sn:0
  //: /line:"26"
  //: /end
  assign Sa = {w52, w96, w240, w234, w228, w92, w91, w195, w89, w159, w216, w86, w204, w84, w192, w82, w81, w174, w168, w78, w156, w76, w75, w74, w73, w136, w71, w124, w126, w120, w67, w66}; //: CONCAT g5  @(1033,1135) /sn:0 /w:[ 5 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:1 /tp:0 /drp:1
  //: joint g79 (C) @(716, 1236) /w:[ -1 26 100 25 ]
  _GGOR2 #(6) g95 (.I0(w32), .I1(w80), .Z(w41));   //: @(303,2415) /sn:0 /w:[ 5 7 0 ]
  //: comment g117 @(350,27) /sn:0
  //: /line:"4"
  //: /end
  ALU1bit g36 (.C(C), .AcarreoE(w173), .B(w178), .A(w16), .AcarreoS(w179), .Sa(w81));   //: @(370, 1000) /sz:(87, 60) /sn:0 /p:[ Ti0>95 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  ALU1bit g24 (.AcarreoE(w122), .C(C), .A(w4), .B(w36), .AcarreoS(w125), .Sa(w126));   //: @(367, -62) /sz:(87, 60) /sn:0 /p:[ Ti0>1 Ti1>71 Li0>1 Li1>0 Bo0<0 Ro0<1 ]
  //: joint g85 (C) @(716, 1746) /w:[ -1 14 112 13 ]
  Suma g92 (.AcarreoE(w245), .A(w32), .B(w55), .AcarreoS(w59), .Suma(w65));   //: @(333, 2466) /sz:(67, 60) /sn:0 /p:[ Ti0>1 Li0>0 Li1>1 Bo0<0 Ro0<9 ]
  //: joint g144 (w49) @(439, 2432) /w:[ 1 2 -1 4 ]
  //: comment g125 @(380,735) /sn:0
  //: /line:"12"
  //: /end
  //: comment g60 @(360,1587) /sn:0
  //: /line:"22"
  //: /end
  //: joint g81 (C) @(716, 1414) /w:[ -1 22 104 21 ]
  _GGNBUF #(2) g101 (.I(w80), .Z(w68));   //: @(163,2556) /sn:0 /w:[ 15 0 ]
  ALU1bit g45 (.C(C), .AcarreoE(w175), .B(w57), .A(w25), .AcarreoS(w193), .Sa(w195));   //: @(385, 1754) /sz:(87, 60) /sn:0 /p:[ Ti0>113 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<0 ]
  //: comment g126 @(375,809) /sn:0
  //: /line:"13"
  //: /end
  //: joint g70 (C) @(716, 459) /w:[ -1 44 82 43 ]
  //: joint g22 (w33) @(228, -324) /w:[ 6 -1 5 8 ]
  ALU1bit g35 (.C(C), .AcarreoE(w167), .B(w172), .A(w15), .AcarreoS(w173), .Sa(w174));   //: @(374, 914) /sz:(87, 60) /sn:0 /p:[ Ti0>93 Ti1>0 Li0>1 Li1>0 Bo0<1 Ro0<1 ]
  //: comment g120 @(356,294) /sn:0
  //: /line:"7"
  //: /end
  //: comment g114 @(353,-261) /sn:0
  //: /line:"1"
  //: /end
  //: GROUND g97 (w49) @(451,2504) /sn:0 /w:[ 13 ]
  //: joint g66 (C) @(717, 104) /w:[ -1 52 74 51 ]
  //: joint g12 (w33) @(305, -376) /w:[ 1 -1 2 12 ]
  //: joint g18 (w2) @(530, -464) /w:[ -1 4 3 6 ]
  //: OUT g108 (Overflow) @(410,2708) /sn:0 /w:[ 1 ]
  ALU1bit g30 (.C(C), .AcarreoE(w141), .B(w152), .A(w9), .AcarreoS(w143), .Sa(w74));   //: @(372, 394) /sz:(87, 60) /sn:0 /p:[ Ti0>81 Ti1>1 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  //: comment g118 @(351,115) /sn:0
  //: /line:"5"
  //: /end
  //: comment g134 @(371,1496) /sn:0
  //: /line:"21"
  //: /end

endmodule
//: /netlistEnd

//: /netlistBegin Mux3x5
module Mux3x5(E0, C, E1, E6, E2, E4, E7, Sa, E5, E3);
//: interface  /sz:(40, 160) /bd:[ Ti0>C[2:0](20/40) Li0>E0[4:0](16/160) Li1>E1[4:0](32/160) Li2>E2[4:0](48/160) Li3>E3[4:0](64/160) Li4>E4[4:0](87/160) Li5>E5[4:0](104/160) Li6>E6[4:0](122/160) Li7>E7[4:0](143/160) Ro0<Sa[4:0](99/160) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [4:0] E7;    //: /sn:0 {0}(#:-103,948)(-88,948)(-88,951)(#:-51,951){1}
input [4:0] E1;    //: /sn:0 {0}(#:42,-154)(92,-154)(92,-157)(#:105,-157){1}
supply0 w0;    //: /sn:0 {0}(213,-303)(193,-303)(193,-305)(183,-305){1}
//: {2}(181,-307)(181,-323)(213,-323){3}
//: {4}(183,-305)(173,-305)(173,-313)(213,-313){5}
//: {6}(181,-303)(181,-287){7}
//: {8}(183,-285)(193,-285)(193,-283)(213,-283){9}
//: {10}(179,-285)(169,-285)(169,-293)(213,-293){11}
//: {12}(181,-283)(181,-265){13}
//: {14}(183,-263)(213,-263){15}
//: {16}(179,-263)(169,-263)(169,-273)(213,-273){17}
//: {18}(181,-261)(181,-247){19}
//: {20}(183,-245)(193,-245)(193,-243)(213,-243){21}
//: {22}(179,-245)(169,-245)(169,-253)(213,-253){23}
//: {24}(181,-243)(181,-225){25}
//: {26}(183,-223)(213,-223){27}
//: {28}(179,-223)(169,-223)(169,-233)(213,-233){29}
//: {30}(181,-221)(181,-205){31}
//: {32}(183,-203)(213,-203){33}
//: {34}(179,-203)(169,-203)(169,-213)(213,-213){35}
//: {36}(181,-201)(181,-188){37}
//: {38}(183,-186)(193,-186)(193,-183)(213,-183){39}
//: {40}(183,-186)(173,-186)(173,-193)(213,-193){41}
//: {42}(181,-184)(181,-165){43}
//: {44}(183,-163)(213,-163){45}
//: {46}(183,-163)(173,-163)(173,-173)(213,-173){47}
//: {48}(181,-161)(181,-144){49}
//: {50}(183,-142)(193,-142)(193,-143)(213,-143){51}
//: {52}(183,-142)(173,-142)(173,-153)(213,-153){53}
//: {54}(181,-140)(181,-126){55}
//: {56}(183,-124)(193,-124)(193,-123)(213,-123){57}
//: {58}(183,-124)(173,-124)(173,-133)(213,-133){59}
//: {60}(181,-122)(181,-105){61}
//: {62}(183,-103)(213,-103){63}
//: {64}(183,-103)(173,-103)(173,-113)(213,-113){65}
//: {66}(181,-101)(181,-85){67}
//: {68}(183,-83)(213,-83){69}
//: {70}(179,-83)(169,-83)(169,-93)(213,-93){71}
//: {72}(181,-81)(181,-65){73}
//: {74}(183,-63)(213,-63){75}
//: {76}(179,-63)(171,-63)(171,215)(99,215){77}
//: {78}(97,213)(97,135){79}
//: {80}(99,133)(112,133){81}
//: {82}(116,133)(151,133){83}
//: {84}(114,131)(114,115){85}
//: {86}(116,113)(151,113){87}
//: {88}(114,111)(114,95){89}
//: {90}(116,93)(151,93){91}
//: {92}(114,91)(114,74){93}
//: {94}(116,72)(126,72)(126,73)(151,73){95}
//: {96}(114,70)(114,52){97}
//: {98}(116,50)(126,50)(126,53)(151,53){99}
//: {100}(114,48)(114,24){101}
//: {102}(116,22)(126,22)(126,23)(151,23){103}
//: {104}(114,20)(114,1){105}
//: {106}(116,-1)(126,-1)(126,3)(151,3){107}
//: {108}(114,-3)(114,-18){109}
//: {110}(116,-20)(126,-20)(126,-17)(151,-17){111}
//: {112}(114,-22)(114,-34){113}
//: {114}(116,-36)(126,-36)(126,-37)(151,-37){115}
//: {116}(114,-38)(114,-48){117}
//: {118}(116,-50)(126,-50)(126,-47)(151,-47){119}
//: {120}(114,-52)(114,-77){121}
//: {122}(116,-79)(126,-79)(126,-77)(151,-77){123}
//: {124}(114,-81)(114,-96){125}
//: {126}(116,-98)(126,-98)(126,-97)(151,-97){127}
//: {128}(114,-100)(114,-114){129}
//: {130}(116,-116)(126,-116)(126,-117)(151,-117){131}
//: {132}(114,-118)(114,-127)(151,-127){133}
//: {134}(116,-116)(106,-116)(106,-107)(151,-107){135}
//: {136}(116,-98)(106,-98)(106,-87)(151,-87){137}
//: {138}(116,-79)(106,-79)(106,-67)(151,-67){139}
//: {140}(112,-50)(102,-50)(102,-57)(151,-57){141}
//: {142}(112,-36)(102,-36)(102,-27)(151,-27){143}
//: {144}(116,-20)(106,-20)(106,-7)(151,-7){145}
//: {146}(116,-1)(106,-1)(106,13)(151,13){147}
//: {148}(116,22)(106,22)(106,33)(151,33){149}
//: {150}(116,50)(106,50)(106,43)(151,43){151}
//: {152}(112,72)(101,72)(101,83)(151,83){153}
//: {154}(116,93)(106,93)(106,103)(151,103){155}
//: {156}(116,113)(106,113)(106,123)(151,123){157}
//: {158}(97,131)(97,63)(151,63){159}
//: {160}(97,217)(97,363)(24,363){161}
//: {162}(22,361)(22,302){163}
//: {164}(24,300)(34,300)(34,302)(73,302){165}
//: {166}(22,298)(22,283){167}
//: {168}(24,281)(34,281)(34,282)(73,282){169}
//: {170}(22,279)(22,264){171}
//: {172}(24,262)(73,262){173}
//: {174}(22,260)(22,244){175}
//: {176}(24,242)(73,242){177}
//: {178}(22,240)(22,224){179}
//: {180}(24,222)(73,222){181}
//: {182}(22,220)(22,204){183}
//: {184}(24,202)(73,202){185}
//: {186}(22,200)(22,183){187}
//: {188}(24,181)(34,181)(34,182)(73,182){189}
//: {190}(22,179)(22,164){191}
//: {192}(24,162)(73,162){193}
//: {194}(22,160)(22,143){195}
//: {196}(24,141)(34,141)(34,142)(73,142){197}
//: {198}(22,139)(22,122){199}
//: {200}(24,120)(34,120)(34,122)(73,122){201}
//: {202}(22,118)(22,104){203}
//: {204}(24,102)(73,102){205}
//: {206}(22,100)(22,83){207}
//: {208}(24,81)(34,81)(34,82)(73,82){209}
//: {210}(22,79)(22,64){211}
//: {212}(24,62)(73,62){213}
//: {214}(22,60)(22,42)(73,42){215}
//: {216}(24,62)(14,62)(14,52)(73,52){217}
//: {218}(24,81)(14,81)(14,72)(73,72){219}
//: {220}(24,102)(14,102)(14,92)(73,92){221}
//: {222}(24,120)(14,120)(14,112)(73,112){223}
//: {224}(24,141)(14,141)(14,132)(73,132){225}
//: {226}(24,162)(14,162)(14,152)(73,152){227}
//: {228}(20,181)(10,181)(10,172)(73,172){229}
//: {230}(24,202)(14,202)(14,192)(73,192){231}
//: {232}(24,222)(14,222)(14,212)(73,212){233}
//: {234}(24,242)(14,242)(14,232)(73,232){235}
//: {236}(24,262)(14,262)(14,252)(73,252){237}
//: {238}(24,281)(14,281)(14,272)(73,272){239}
//: {240}(24,300)(14,300)(14,292)(73,292){241}
//: {242}(22,365)(22,509){243}
//: {244}(24,511)(90,511)(90,469)(107,469){245}
//: {246}(111,469)(152,469){247}
//: {248}(156,469)(170,469)(170,468)(184,468){249}
//: {250}(154,467)(154,452){251}
//: {252}(156,450)(178,450)(178,448)(184,448){253}
//: {254}(154,448)(154,431){255}
//: {256}(156,429)(170,429)(170,428)(184,428){257}
//: {258}(154,427)(154,411){259}
//: {260}(156,409)(172,409)(172,408)(184,408){261}
//: {262}(154,407)(154,391){263}
//: {264}(156,389)(170,389)(170,388)(184,388){265}
//: {266}(154,387)(154,372){267}
//: {268}(156,370)(170,370)(170,368)(184,368){269}
//: {270}(154,368)(154,353){271}
//: {272}(156,351)(172,351)(172,348)(184,348){273}
//: {274}(154,349)(154,338)(184,338){275}
//: {276}(152,351)(146,351)(146,358)(184,358){277}
//: {278}(152,370)(146,370)(146,378)(184,378){279}
//: {280}(152,389)(146,389)(146,398)(184,398){281}
//: {282}(152,409)(146,409)(146,418)(184,418){283}
//: {284}(152,429)(146,429)(146,438)(184,438){285}
//: {286}(152,450)(142,450)(142,458)(184,458){287}
//: {288}(154,471)(154,485){289}
//: {290}(156,487)(166,487)(166,488)(184,488){291}
//: {292}(152,487)(142,487)(142,498)(184,498){293}
//: {294}(154,489)(154,506){295}
//: {296}(156,508)(184,508){297}
//: {298}(152,508)(142,508)(142,518)(184,518){299}
//: {300}(154,510)(154,526){301}
//: {302}(156,528)(184,528){303}
//: {304}(152,528)(142,528)(142,538)(184,538){305}
//: {306}(154,530)(154,545){307}
//: {308}(156,547)(166,547)(166,548)(184,548){309}
//: {310}(156,547)(146,547)(146,558)(184,558){311}
//: {312}(154,549)(154,564){313}
//: {314}(156,566)(166,566)(166,568)(184,568){315}
//: {316}(156,566)(146,566)(146,578)(184,578){317}
//: {318}(154,568)(154,599){319}
//: {320}(156,601)(172,601)(172,598)(184,598){321}
//: {322}(156,601)(146,601)(146,588)(184,588){323}
//: {324}(154,603)(154,861)(82,861){325}
//: {326}(80,859)(80,842)(84,842){327}
//: {328}(88,842)(96,842)(96,841)(123,841){329}
//: {330}(86,840)(86,831)(123,831){331}
//: {332}(86,844)(86,850)(105,850)(105,834)(89,834)(89,822){333}
//: {334}(91,820)(101,820)(101,821)(123,821){335}
//: {336}(89,818)(89,803){337}
//: {338}(91,801)(123,801){339}
//: {340}(89,799)(89,781){341}
//: {342}(91,779)(101,779)(101,781)(123,781){343}
//: {344}(89,777)(89,762){345}
//: {346}(91,760)(101,760)(101,761)(123,761){347}
//: {348}(89,758)(89,743){349}
//: {350}(91,741)(123,741){351}
//: {352}(89,739)(89,723){353}
//: {354}(91,721)(123,721){355}
//: {356}(89,719)(89,691){357}
//: {358}(91,689)(101,689)(101,691)(123,691){359}
//: {360}(89,687)(89,672){361}
//: {362}(91,670)(101,670)(101,671)(123,671){363}
//: {364}(89,668)(89,651){365}
//: {366}(91,649)(101,649)(101,651)(123,651){367}
//: {368}(89,647)(89,631){369}
//: {370}(91,629)(101,629)(101,631)(123,631){371}
//: {372}(89,627)(89,612){373}
//: {374}(91,610)(101,610)(101,611)(123,611){375}
//: {376}(89,608)(89,591)(103,591){377}
//: {378}(107,591)(123,591){379}
//: {380}(105,589)(105,581)(123,581){381}
//: {382}(105,593)(105,601)(123,601){383}
//: {384}(91,610)(81,610)(81,621)(123,621){385}
//: {386}(87,629)(76,629)(76,641)(123,641){387}
//: {388}(91,649)(81,649)(81,661)(123,661){389}
//: {390}(91,670)(81,670)(81,681)(123,681){391}
//: {392}(91,689)(81,689)(81,701)(123,701){393}
//: {394}(87,721)(77,721)(77,711)(123,711){395}
//: {396}(91,741)(81,741)(81,731)(123,731){397}
//: {398}(91,760)(81,760)(81,751)(123,751){399}
//: {400}(91,779)(81,779)(81,771)(123,771){401}
//: {402}(91,801)(81,801)(81,791)(123,791){403}
//: {404}(87,820)(77,820)(77,811)(123,811){405}
//: {406}(80,863)(80,1047)(33,1047){407}
//: {408}(31,1045)(31,1027){409}
//: {410}(33,1025)(64,1025){411}
//: {412}(31,1023)(31,1005){413}
//: {414}(33,1003)(42,1003)(42,1005)(64,1005){415}
//: {416}(31,1001)(31,972){417}
//: {418}(33,970)(42,970)(42,975)(64,975){419}
//: {420}(31,968)(31,954){421}
//: {422}(33,952)(42,952)(42,955)(64,955){423}
//: {424}(31,950)(31,938){425}
//: {426}(33,936)(42,936)(42,935)(64,935){427}
//: {428}(31,934)(31,916){429}
//: {430}(33,914)(42,914)(42,915)(64,915){431}
//: {432}(31,912)(31,896){433}
//: {434}(33,894)(42,894)(42,895)(64,895){435}
//: {436}(31,892)(31,877){437}
//: {438}(33,875)(64,875){439}
//: {440}(31,873)(31,856){441}
//: {442}(33,854)(42,854)(42,855)(64,855){443}
//: {444}(31,852)(31,837){445}
//: {446}(33,835)(64,835){447}
//: {448}(31,833)(31,824){449}
//: {450}(33,822)(42,822)(42,825)(64,825){451}
//: {452}(31,820)(31,796){453}
//: {454}(33,794)(42,794)(42,795)(64,795){455}
//: {456}(31,792)(31,778){457}
//: {458}(33,776)(42,776)(42,775)(64,775){459}
//: {460}(31,774)(31,765)(64,765){461}
//: {462}(29,776)(18,776)(18,785)(64,785){463}
//: {464}(29,794)(18,794)(18,805)(64,805){465}
//: {466}(29,822)(18,822)(18,815)(64,815){467}
//: {468}(29,835)(18,835)(18,845)(64,845){469}
//: {470}(29,854)(18,854)(18,865)(64,865){471}
//: {472}(29,875)(18,875)(18,885)(64,885){473}
//: {474}(29,894)(18,894)(18,905)(64,905){475}
//: {476}(29,914)(18,914)(18,925)(64,925){477}
//: {478}(29,936)(18,936)(18,945)(64,945){479}
//: {480}(29,952)(18,952)(18,965)(64,965){481}
//: {482}(29,970)(18,970)(18,985)(64,985){483}
//: {484}(29,1003)(18,1003)(18,988)(46,988)(46,995)(64,995){485}
//: {486}(29,1025)(18,1025)(18,1015)(64,1015){487}
//: {488}(31,1049)(31,1257)(-22,1257){489}
//: {490}(-24,1255)(-24,1241){491}
//: {492}(-22,1239)(-12,1239)(-12,1240)(4,1240){493}
//: {494}(-24,1237)(-24,1208){495}
//: {496}(-22,1206)(-12,1206)(-12,1210)(4,1210){497}
//: {498}(-24,1204)(-24,1190){499}
//: {500}(-22,1188)(-12,1188)(-12,1190)(4,1190){501}
//: {502}(-24,1186)(-24,1171){503}
//: {504}(-22,1169)(-12,1169)(-12,1170)(4,1170){505}
//: {506}(-24,1167)(-24,1151){507}
//: {508}(-22,1149)(-12,1149)(-12,1150)(4,1150){509}
//: {510}(-24,1147)(-24,1131){511}
//: {512}(-22,1129)(-12,1129)(-12,1130)(4,1130){513}
//: {514}(-24,1127)(-24,1110){515}
//: {516}(-22,1108)(-12,1108)(-12,1110)(4,1110){517}
//: {518}(-24,1106)(-24,1092){519}
//: {520}(-22,1090)(4,1090){521}
//: {522}(-24,1088)(-24,1072){523}
//: {524}(-22,1070)(4,1070){525}
//: {526}(-24,1068)(-24,1054){527}
//: {528}(-22,1052)(-12,1052)(-12,1050)(4,1050){529}
//: {530}(-24,1050)(-24,1029){531}
//: {532}(-22,1027)(-12,1027)(-12,1030)(4,1030){533}
//: {534}(-24,1025)(-24,1012){535}
//: {536}(-22,1010)(4,1010){537}
//: {538}(-24,1008)(-24,991){539}
//: {540}(-22,989)(-12,989)(-12,990)(4,990){541}
//: {542}(-24,987)(-24,980)(4,980){543}
//: {544}(-22,989)(-32,989)(-32,1000)(4,1000){545}
//: {546}(-26,1010)(-36,1010)(-36,1020)(4,1020){547}
//: {548}(-26,1027)(-36,1027)(-36,1040)(4,1040){549}
//: {550}(-22,1052)(-32,1052)(-32,1060)(4,1060){551}
//: {552}(-26,1070)(-36,1070)(-36,1080)(4,1080){553}
//: {554}(-22,1090)(-32,1090)(-32,1100)(4,1100){555}
//: {556}(-22,1108)(-32,1108)(-32,1120)(4,1120){557}
//: {558}(-22,1129)(-32,1129)(-32,1140)(4,1140){559}
//: {560}(-22,1149)(-32,1149)(-32,1160)(4,1160){561}
//: {562}(-26,1169)(-36,1169)(-36,1180)(4,1180){563}
//: {564}(-22,1188)(-32,1188)(-32,1200)(4,1200){565}
//: {566}(-22,1206)(-32,1206)(-32,1220)(4,1220){567}
//: {568}(-26,1239)(-36,1239)(-36,1230)(4,1230){569}
//: {570}(-24,1259)(-24,1299){571}
//: {572}(109,471)(109,478)(184,478){573}
//: {574}(20,511)(-99,511)(-99,494)(-70,494){575}
//: {576}(-66,494)(-50,494)(-50,492)(-29,492){577}
//: {578}(-68,492)(-68,482)(-29,482){579}
//: {580}(-68,496)(-68,508)(-82,508)(-82,475){581}
//: {582}(-80,473)(-70,473)(-70,472)(-29,472){583}
//: {584}(-82,471)(-82,454){585}
//: {586}(-80,452)(-29,452){587}
//: {588}(-82,450)(-82,434){589}
//: {590}(-80,432)(-29,432){591}
//: {592}(-82,430)(-82,414){593}
//: {594}(-80,412)(-29,412){595}
//: {596}(-82,410)(-82,384){597}
//: {598}(-80,382)(-29,382){599}
//: {600}(-82,380)(-82,362){601}
//: {602}(-80,360)(-70,360)(-70,362)(-29,362){603}
//: {604}(-82,358)(-82,337){605}
//: {606}(-80,335)(-70,335)(-70,372)(-29,372){607}
//: {608}(-82,333)(-82,323){609}
//: {610}(-80,321)(-70,321)(-70,322)(-29,322){611}
//: {612}(-82,319)(-82,303){613}
//: {614}(-80,301)(-70,301)(-70,302)(-29,302){615}
//: {616}(-82,299)(-82,282){617}
//: {618}(-80,280)(-70,280)(-70,282)(-29,282){619}
//: {620}(-82,278)(-82,261){621}
//: {622}(-80,259)(-70,259)(-70,262)(-29,262){623}
//: {624}(-82,257)(-82,243)(-62,243)(-62,232)(-29,232){625}
//: {626}(-84,259)(-96,259)(-96,252)(-57,252){627}
//: {628}(-53,252)(-29,252){629}
//: {630}(-55,250)(-55,242)(-29,242){631}
//: {632}(-84,280)(-94,280)(-94,272)(-29,272){633}
//: {634}(-80,301)(-90,301)(-90,292)(-29,292){635}
//: {636}(-80,321)(-90,321)(-90,312)(-29,312){637}
//: {638}(-84,335)(-96,335)(-96,342)(-61,342){639}
//: {640}(-57,342)(-29,342){641}
//: {642}(-59,340)(-59,332)(-29,332){643}
//: {644}(-80,360)(-90,360)(-90,352)(-29,352){645}
//: {646}(-84,382)(-94,382)(-94,392)(-29,392){647}
//: {648}(-80,412)(-90,412)(-90,402)(-29,402){649}
//: {650}(-80,432)(-90,432)(-90,422)(-29,422){651}
//: {652}(-80,452)(-90,452)(-90,442)(-29,442){653}
//: {654}(-80,473)(-90,473)(-90,462)(-29,462){655}
//: {656}(181,-61)(181,-51)(196,-51)(196,-73)(213,-73){657}
input [4:0] E2;    //: /sn:0 {0}(#:-42,12)(-13,12)(-13,11)(#:2,11){1}
input [4:0] E0;    //: /sn:0 {0}(#:89,-355)(151,-355)(151,-353)(#:166,-353){1}
input [4:0] E4;    //: /sn:0 {0}(#:70,375)(107,375)(107,310)(#:122,310){1}
output [4:0] Sa;    //: /sn:0 {0}(595,35)(530,35)(#:530,44)(#:515,44){1}
input [2:0] C;    //: /sn:0 {0}(#:324,5)(324,67)(316,67)(#:316,82){1}
input [4:0] E3;    //: /sn:0 {0}(#:-130,212)(-91,212)(-91,202)(#:-76,202){1}
input [4:0] E5;    //: /sn:0 {0}(#:31,567)(59,567)(59,551)(#:74,551){1}
input [4:0] E6;    //: /sn:0 {0}(#:-23,731)(-16,731)(-16,734)(#:9,734){1}
wire [31:0] w6;    //: /sn:0 {0}(#:306,237)(213,237)(213,686)(#:129,686){1}
wire w270;    //: /sn:0 {0}(128,290)(169,290)(169,288)(184,288){1}
wire [31:0] w7;    //: /sn:0 {0}(#:70,870)(220,870)(220,264)(#:306,264){1}
wire w160;    //: /sn:0 {0}(442,201)(457,201){1}
wire w336;    //: /sn:0 {0}(64,715)(38,715)(38,714)(15,714){1}
wire w175;    //: /sn:0 {0}(111,-167)(151,-167){1}
wire w112;    //: /sn:0 {0}(172,-343)(213,-343){1}
wire w166;    //: /sn:0 {0}(442,261)(457,261){1}
wire w339;    //: /sn:0 {0}(15,744)(49,744)(49,745)(64,745){1}
wire w141;    //: /sn:0 {0}(8,-9)(62,-9)(62,-8)(73,-8){1}
wire w153;    //: /sn:0 {0}(442,131)(457,131){1}
wire [31:0] w4;    //: /sn:0 {0}(#:-23,337)(88,337)(88,174)(#:306,174){1}
wire w306;    //: /sn:0 {0}(80,561)(123,561){1}
wire w109;    //: /sn:0 {0}(172,-373)(213,-373){1}
wire w152;    //: /sn:0 {0}(442,121)(457,121){1}
wire w304;    //: /sn:0 {0}(80,541)(123,541){1}
wire w239;    //: /sn:0 {0}(-70,202)(-29,202){1}
wire w207;    //: /sn:0 {0}(8,11)(58,11)(58,12)(73,12){1}
wire w373;    //: /sn:0 {0}(-45,971)(-11,971)(-11,970)(4,970){1}
wire [31:0] w3;    //: /sn:0 {0}(#:79,147)(170,147)(170,148)(#:306,148){1}
wire w151;    //: /sn:0 {0}(442,111)(457,111){1}
wire w271;    //: /sn:0 {0}(128,300)(169,300)(169,298)(184,298){1}
wire w177;    //: /sn:0 {0}(151,-147)(111,-147){1}
wire w240;    //: /sn:0 {0}(-70,212)(-29,212){1}
wire w159;    //: /sn:0 {0}(442,191)(457,191){1}
wire w171;    //: /sn:0 {0}(442,311)(457,311){1}
wire w168;    //: /sn:0 {0}(442,281)(457,281){1}
wire w111;    //: /sn:0 {0}(172,-353)(213,-353){1}
wire w340;    //: /sn:0 {0}(64,755)(29,755)(29,754)(15,754){1}
wire w157;    //: /sn:0 {0}(442,171)(457,171){1}
wire w237;    //: /sn:0 {0}(-70,182)(-29,182){1}
wire w170;    //: /sn:0 {0}(442,301)(457,301){1}
wire w209;    //: /sn:0 {0}(8,31)(58,31)(58,32)(73,32){1}
wire w176;    //: /sn:0 {0}(111,-157)(151,-157){1}
wire w156;    //: /sn:0 {0}(442,161)(457,161){1}
wire w307;    //: /sn:0 {0}(80,571)(123,571){1}
wire w169;    //: /sn:0 {0}(442,291)(457,291){1}
wire w167;    //: /sn:0 {0}(442,271)(457,271){1}
wire w174;    //: /sn:0 {0}(111,-177)(151,-177){1}
wire w161;    //: /sn:0 {0}(442,211)(457,211){1}
wire [31:0] w1;    //: /sn:0 {0}(#:219,-218)(293,-218)(293,106)(#:306,106){1}
wire w241;    //: /sn:0 {0}(-70,222)(-29,222){1}
wire w272;    //: /sn:0 {0}(128,310)(169,310)(169,308)(184,308){1}
wire w369;    //: /sn:0 {0}(-45,931)(-11,931)(-11,930)(4,930){1}
wire w154;    //: /sn:0 {0}(442,141)(457,141){1}
wire w372;    //: /sn:0 {0}(4,960)(-30,960)(-30,961)(-45,961){1}
wire w303;    //: /sn:0 {0}(80,531)(123,531){1}
wire w158;    //: /sn:0 {0}(442,181)(457,181){1}
wire [31:0] w8;    //: /sn:0 {0}(#:10,1085)(291,1085)(291,292)(#:306,292){1}
wire w338;    //: /sn:0 {0}(64,735)(29,735)(29,734)(15,734){1}
wire w164;    //: /sn:0 {0}(442,241)(457,241){1}
wire w371;    //: /sn:0 {0}(-45,951)(-11,951)(-11,950)(4,950){1}
wire w163;    //: /sn:0 {0}(442,231)(457,231){1}
wire w162;    //: /sn:0 {0}(442,221)(457,221){1}
wire w238;    //: /sn:0 {0}(-70,192)(-29,192){1}
wire w144;    //: /sn:0 {0}(509,44)(457,44)(457,41)(442,41){1}
wire w149;    //: /sn:0 {0}(442,91)(457,91){1}
wire w146;    //: /sn:0 {0}(442,61)(496,61)(496,64)(509,64){1}
wire w165;    //: /sn:0 {0}(442,251)(457,251){1}
wire w172;    //: /sn:0 {0}(442,321)(457,321){1}
wire w173;    //: /sn:0 {0}(442,331)(457,331){1}
wire [31:0] w2;    //: /sn:0 {0}(#:157,-22)(253,-22)(253,126)(#:306,126){1}
wire w113;    //: /sn:0 {0}(172,-333)(213,-333){1}
wire w150;    //: /sn:0 {0}(442,101)(457,101){1}
wire w110;    //: /sn:0 {0}(172,-363)(213,-363){1}
wire w148;    //: /sn:0 {0}(442,81)(457,81){1}
wire w206;    //: /sn:0 {0}(8,1)(58,1)(58,2)(73,2){1}
wire w274;    //: /sn:0 {0}(128,330)(169,330)(169,328)(184,328){1}
wire w273;    //: /sn:0 {0}(128,320)(169,320)(169,318)(184,318){1}
wire w208;    //: /sn:0 {0}(8,21)(58,21)(58,22)(73,22){1}
wire [31:0] w5;    //: /sn:0 {0}(#:190,443)(196,443)(196,212)(#:306,212){1}
wire w143;    //: /sn:0 {0}(509,34)(457,34)(457,31)(442,31){1}
wire w178;    //: /sn:0 {0}(111,-137)(151,-137){1}
wire w155;    //: /sn:0 {0}(442,151)(457,151){1}
wire w142;    //: /sn:0 {0}(509,24)(457,24)(457,21)(442,21){1}
wire w147;    //: /sn:0 {0}(442,71)(457,71){1}
wire w145;    //: /sn:0 {0}(509,54)(457,54)(457,51)(442,51){1}
wire [31:0] w9;    //: /sn:0 {0}(#:348,176)(#:436,176){1}
wire w370;    //: /sn:0 {0}(4,940)(-30,940)(-30,941)(-45,941){1}
wire w337;    //: /sn:0 {0}(15,724)(49,724)(49,725)(64,725){1}
wire w305;    //: /sn:0 {0}(80,551)(123,551){1}
//: enddecls

  assign w1 = {w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w113, w112, w111, w110, w109}; //: CONCAT g4  @(218,-218) /sn:0 /w:[ 0 75 657 69 71 63 65 57 59 51 53 45 47 39 41 33 35 27 29 21 23 15 17 9 11 0 5 3 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign w4 = {w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w241, w240, w239, w238, w237}; //: CONCAT g8  @(-24,337) /sn:0 /w:[ 0 577 579 583 655 587 653 591 651 595 649 647 599 607 603 645 641 643 611 637 615 635 619 633 623 629 631 625 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: joint g140 (w0) @(181, -285) /w:[ 8 7 10 12 ]
  assign {w209, w208, w207, w206, w141} = E2; //: CONCAT g13  @(3,11) /sn:0 /R:2 /w:[ 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: joint g37 (w0) @(-24, 1169) /w:[ 504 506 562 503 ]
  //: joint g55 (w0) @(31, 1047) /w:[ 407 408 -1 488 ]
  //: joint g58 (w0) @(89, 820) /w:[ 334 336 404 333 ]
  //: joint g139 (w0) @(181, -263) /w:[ 14 13 16 18 ]
  assign Sa = {w146, w145, w144, w143, w142}; //: CONCAT g112  @(514,44) /sn:0 /w:[ 1 1 0 0 0 0 ] /dr:1 /tp:0 /drp:1
  //: joint g76 (w0) @(154, 450) /w:[ 252 254 286 251 ]
  //: joint g111 (w0) @(22, 62) /w:[ 212 214 216 211 ]
  assign w2 = {w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w178, w177, w176, w175, w174}; //: CONCAT g1  @(156,-22) /sn:0 /w:[ 0 83 157 87 155 91 153 95 159 99 151 149 103 147 107 145 111 143 115 119 141 139 123 137 127 135 131 133 1 0 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: joint g64 (w0) @(89, 610) /w:[ 374 376 384 373 ]
  assign w7 = {w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w340, w339, w338, w337, w336}; //: CONCAT g11  @(69,870) /sn:0 /w:[ 0 411 487 415 485 483 419 481 423 479 427 477 431 475 435 473 439 471 443 469 447 451 467 465 455 463 459 461 0 1 0 1 0 ] /dr:1 /tp:0 /drp:1
  //: joint g130 (w0) @(181, -83) /w:[ 68 67 70 72 ]
  //: joint g121 (w0) @(114, -79) /w:[ 122 124 138 121 ]
  //: joint g28 (w0) @(-24, 989) /w:[ 540 542 544 539 ]
  //: joint g50 (w0) @(31, 914) /w:[ 430 432 476 429 ]
  //: joint g132 (w0) @(181, -124) /w:[ 56 55 58 60 ]
  //: IN g19 (E0) @(87,-355) /sn:0 /w:[ 0 ]
  //: joint g113 (w0) @(22, 363) /w:[ 161 162 -1 242 ]
  //: IN g6 (C) @(324,3) /sn:0 /R:3 /w:[ 0 ]
  //: joint g38 (w0) @(-24, 1188) /w:[ 500 502 564 499 ]
  //: joint g115 (w0) @(114, 113) /w:[ 86 88 156 85 ]
  assign {w178, w177, w176, w175, w174} = E1; //: CONCAT g7  @(106,-157) /sn:0 /R:2 /w:[ 0 1 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: joint g53 (w0) @(31, 970) /w:[ 418 420 482 417 ]
  //: joint g75 (w0) @(154, 429) /w:[ 256 258 284 255 ]
  //: joint g135 (w0) @(181, -186) /w:[ 38 37 40 42 ]
  //: IN g20 (E1) @(40,-154) /sn:0 /w:[ 0 ]
  //: joint g31 (w0) @(-24, 1052) /w:[ 528 530 550 527 ]
  //: joint g124 (w0) @(114, -20) /w:[ 110 112 144 109 ]
  //: joint g39 (w0) @(-24, 1206) /w:[ 496 498 566 495 ]
  //: joint g68 (w0) @(89, 689) /w:[ 358 360 392 357 ]
  //: joint g48 (w0) @(31, 875) /w:[ 438 440 472 437 ]
  assign {w340, w339, w338, w337, w336} = E6; //: CONCAT g17  @(10,734) /sn:0 /R:2 /w:[ 1 0 1 0 1 1 ] /dr:0 /tp:0 /drp:0
  //: IN g25 (E6) @(-25,731) /sn:0 /w:[ 0 ]
  //: joint g29 (w0) @(-24, 1010) /w:[ 536 538 546 535 ]
  //: joint g52 (w0) @(31, 952) /w:[ 422 424 480 421 ]
  //: joint g106 (w0) @(22, 162) /w:[ 192 194 226 191 ]
  //: joint g107 (w0) @(22, 141) /w:[ 196 198 224 195 ]
  //: joint g83 (w0) @(109, 469) /w:[ 246 -1 245 572 ]
  //: joint g100 (w0) @(22, 281) /w:[ 168 170 238 167 ]
  assign {w241, w240, w239, w238, w237} = E3; //: CONCAT g14  @(-75,202) /sn:0 /R:2 /w:[ 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: joint g44 (w0) @(31, 794) /w:[ 454 456 464 453 ]
  //: joint g47 (w0) @(31, 854) /w:[ 442 444 470 441 ]
  //: joint g80 (w0) @(154, 528) /w:[ 302 301 304 306 ]
  //: joint g94 (w0) @(-82, 301) /w:[ 614 616 634 613 ]
  //: IN g21 (E2) @(-44,12) /sn:0 /w:[ 0 ]
  //: joint g84 (w0) @(-68, 494) /w:[ 576 578 575 580 ]
  //: joint g105 (w0) @(22, 181) /w:[ 188 190 228 187 ]
  //: joint g141 (w0) @(181, -305) /w:[ 1 2 4 6 ]
  //: IN g23 (E4) @(68,375) /sn:0 /w:[ 0 ]
  //: joint g41 (w0) @(-24, 1257) /w:[ 489 490 -1 570 ]
  //: joint g40 (w0) @(-24, 1239) /w:[ 492 494 568 491 ]
  //: joint g54 (w0) @(31, 1003) /w:[ 414 416 484 413 ]
  //: joint g93 (w0) @(-82, 321) /w:[ 610 612 636 609 ]
  //: joint g116 (w0) @(114, 93) /w:[ 90 92 154 89 ]
  //: joint g123 (w0) @(114, -36) /w:[ 114 116 142 113 ]
  Mux3x32 g0 (.C(C), .E7(w8), .E6(w7), .E5(w6), .E4(w5), .E3(w4), .E2(w3), .E1(w2), .E0(w1), .Sa(w9));   //: @(307, 83) /sz:(40, 234) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Li2>0 Li3>1 Li4>1 Li5>1 Li6>1 Li7>1 Ro0<0 ]
  //: IN g26 (E7) @(-105,948) /sn:0 /w:[ 0 ]
  //: joint g46 (w0) @(31, 835) /w:[ 446 448 468 445 ]
  //: joint g90 (w0) @(-82, 335) /w:[ 606 608 638 605 ]
  //: joint g82 (w0) @(154, 566) /w:[ 314 313 316 318 ]
  //: joint g136 (w0) @(181, -203) /w:[ 32 31 34 36 ]
  //: joint g128 (w0) @(97, 215) /w:[ 77 78 -1 160 ]
  //: joint g33 (w0) @(-24, 1090) /w:[ 520 522 554 519 ]
  //: joint g91 (w0) @(-82, 360) /w:[ 602 604 644 601 ]
  //: joint g49 (w0) @(31, 894) /w:[ 434 436 474 433 ]
  //: joint g137 (w0) @(181, -223) /w:[ 26 25 28 30 ]
  //: joint g61 (w0) @(89, 760) /w:[ 346 348 398 345 ]
  assign {w113, w112, w111, w110, w109} = E0; //: CONCAT g3  @(167,-353) /sn:0 /R:2 /w:[ 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: joint g34 (w0) @(-24, 1108) /w:[ 516 518 556 515 ]
  //: joint g51 (w0) @(31, 936) /w:[ 426 428 478 425 ]
  //: joint g86 (w0) @(-82, 452) /w:[ 586 588 652 585 ]
  //: joint g89 (w0) @(-82, 382) /w:[ 598 600 646 597 ]
  assign w3 = {w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w209, w208, w207, w206, w141}; //: CONCAT g2  @(78,147) /sn:0 /w:[ 0 165 241 169 239 173 237 177 235 181 233 185 231 189 229 193 227 197 225 201 223 205 221 209 219 213 217 215 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: joint g65 (w0) @(89, 629) /w:[ 370 372 386 369 ]
  //: joint g77 (w0) @(154, 469) /w:[ 248 250 247 288 ]
  //: joint g110 (w0) @(22, 81) /w:[ 208 210 218 207 ]
  //: joint g59 (w0) @(89, 801) /w:[ 338 340 402 337 ]
  //: joint g72 (w0) @(154, 370) /w:[ 268 270 278 267 ]
  //: joint g98 (w0) @(22, 511) /w:[ 244 243 574 -1 ]
  //: joint g99 (w0) @(22, 300) /w:[ 164 166 240 163 ]
  assign {w307, w306, w305, w304, w303} = E5; //: CONCAT g16  @(75,551) /sn:0 /R:2 /w:[ 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: joint g96 (w0) @(-82, 259) /w:[ 622 624 626 621 ]
  //: joint g103 (w0) @(22, 222) /w:[ 180 182 232 179 ]
  //: joint g122 (w0) @(114, -50) /w:[ 118 120 140 117 ]
  assign w6 = {w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w307, w306, w305, w304, w303}; //: CONCAT g10  @(128,686) /sn:0 /w:[ 1 329 331 335 405 339 403 343 401 347 399 351 397 355 395 393 359 391 363 389 367 387 371 385 375 383 379 381 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: joint g78 (w0) @(154, 487) /w:[ 290 289 292 294 ]
  //: joint g87 (w0) @(-82, 432) /w:[ 590 592 650 589 ]
  //: joint g129 (w0) @(181, -63) /w:[ 74 73 76 656 ]
  //: GROUND g27 (w0) @(-24,1305) /sn:0 /w:[ 571 ]
  //: joint g32 (w0) @(-24, 1070) /w:[ 524 526 552 523 ]
  //: joint g102 (w0) @(22, 242) /w:[ 176 178 234 175 ]
  //: joint g69 (w0) @(80, 861) /w:[ 325 326 -1 406 ]
  assign w5 = {w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w274, w273, w272, w271, w270}; //: CONCAT g9  @(189,443) /sn:0 /w:[ 0 321 323 317 315 311 309 305 303 299 297 293 291 573 249 287 253 285 257 283 261 281 265 279 269 277 273 275 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: joint g57 (w0) @(105, 591) /w:[ 378 380 377 382 ]
  //: joint g119 (w0) @(114, -116) /w:[ 130 132 134 129 ]
  //: OUT g142 (Sa) @(592,35) /sn:0 /w:[ 0 ]
  assign {w274, w273, w272, w271, w270} = E4; //: CONCAT g15  @(123,310) /sn:0 /R:2 /w:[ 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: joint g71 (w0) @(154, 351) /w:[ 272 274 276 271 ]
  //: joint g131 (w0) @(181, -103) /w:[ 62 61 64 66 ]
  //: joint g67 (w0) @(89, 670) /w:[ 362 364 390 361 ]
  //: joint g127 (w0) @(97, 133) /w:[ 80 158 -1 79 ]
  //: joint g43 (w0) @(31, 776) /w:[ 458 460 462 457 ]
  //: joint g62 (w0) @(89, 741) /w:[ 350 352 396 349 ]
  //: joint g73 (w0) @(154, 389) /w:[ 264 266 280 263 ]
  //: joint g88 (w0) @(-82, 412) /w:[ 594 596 648 593 ]
  //: joint g104 (w0) @(22, 202) /w:[ 184 186 230 183 ]
  //: joint g138 (w0) @(181, -245) /w:[ 20 19 22 24 ]
  //: joint g42 (w0) @(31, 1025) /w:[ 410 412 486 409 ]
  //: joint g63 (w0) @(89, 721) /w:[ 354 356 394 353 ]
  //: joint g74 (w0) @(154, 409) /w:[ 260 262 282 259 ]
  //: joint g109 (w0) @(22, 102) /w:[ 204 206 220 203 ]
  //: joint g133 (w0) @(181, -142) /w:[ 50 49 52 54 ]
  assign {w173, w172, w171, w170, w169, w168, w167, w166, w165, w164, w163, w162, w161, w160, w159, w158, w157, w156, w155, w154, w153, w152, w151, w150, w149, w148, w147, w146, w145, w144, w143, w142} = w9; //: CONCAT g5  @(437,176) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 ] /dr:0 /tp:0 /drp:0
  //: joint g56 (w0) @(86, 842) /w:[ 328 330 327 332 ]
  //: joint g79 (w0) @(154, 508) /w:[ 296 295 298 300 ]
  //: joint g95 (w0) @(-82, 280) /w:[ 618 620 632 617 ]
  //: joint g117 (w0) @(114, 72) /w:[ 94 96 152 93 ]
  //: IN g24 (E5) @(29,567) /sn:0 /w:[ 0 ]
  //: joint g36 (w0) @(-24, 1149) /w:[ 508 510 560 507 ]
  //: joint g85 (w0) @(-82, 473) /w:[ 582 584 654 581 ]
  //: joint g92 (w0) @(-59, 342) /w:[ 640 642 639 -1 ]
  //: joint g125 (w0) @(114, -1) /w:[ 106 108 146 105 ]
  //: joint g60 (w0) @(89, 779) /w:[ 342 344 400 341 ]
  //: joint g81 (w0) @(154, 547) /w:[ 308 307 310 312 ]
  //: joint g101 (w0) @(22, 262) /w:[ 172 174 236 171 ]
  //: joint g126 (w0) @(114, 22) /w:[ 102 104 148 101 ]
  //: joint g70 (w0) @(154, 601) /w:[ 320 319 322 324 ]
  //: joint g45 (w0) @(31, 822) /w:[ 450 452 466 449 ]
  //: joint g35 (w0) @(-24, 1129) /w:[ 512 514 558 511 ]
  //: IN g22 (E3) @(-132,212) /sn:0 /w:[ 0 ]
  //: joint g120 (w0) @(114, -98) /w:[ 126 128 136 125 ]
  //: joint g114 (w0) @(114, 133) /w:[ 82 84 81 -1 ]
  //: joint g97 (w0) @(-55, 252) /w:[ 628 630 627 -1 ]
  //: joint g66 (w0) @(89, 649) /w:[ 366 368 388 365 ]
  assign {w373, w372, w371, w370, w369} = E7; //: CONCAT g18  @(-50,951) /sn:0 /R:2 /w:[ 0 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  assign w8 = {w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w0, w373, w372, w371, w370, w369}; //: CONCAT g12  @(9,1085) /sn:0 /w:[ 0 493 569 567 497 565 501 563 505 561 509 559 513 557 517 555 521 553 525 551 529 549 533 547 537 545 541 543 1 0 1 0 1 ] /dr:1 /tp:0 /drp:1
  //: joint g108 (w0) @(22, 120) /w:[ 200 202 222 199 ]
  //: joint g30 (w0) @(-24, 1027) /w:[ 532 534 548 531 ]
  //: joint g118 (w0) @(114, 50) /w:[ 98 100 150 97 ]
  //: joint g134 (w0) @(181, -163) /w:[ 44 43 46 48 ]

endmodule
//: /netlistEnd

//: /netlistBegin Extensor16a32
module Extensor16a32(Sa, E);
//: interface  /sz:(97, 40) /bd:[ Li0>E[15:0](16/40) Ro0<Sa[31:0](16/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output [31:0] Sa;    //: /sn:0 {0}(527,346)(463,346)(#:463,257){1}
input [15:0] E;    //: /sn:0 {0}(#:388,124)(543,124)(#:543,197){1}
wire w6;    //: /sn:0 {0}(598,251)(598,203){1}
wire w7;    //: /sn:0 {0}(588,251)(588,203){1}
wire w14;    //: /sn:0 {0}(518,251)(518,203){1}
wire w16;    //: /sn:0 {0}(498,251)(498,203){1}
wire w15;    //: /sn:0 {0}(508,251)(508,203){1}
wire w19;    //: /sn:0 {0}(438,251)(438,236)(437,236)(437,226){1}
//: {2}(439,224)(466,224){3}
//: {4}(470,224)(472,224)(472,232)(458,232)(458,251){5}
//: {6}(468,222)(468,203){7}
//: {8}(468,226)(468,251){9}
//: {10}(437,222)(437,212)(448,212)(448,251){11}
//: {12}(435,224)(419,224){13}
//: {14}(417,222)(417,212)(428,212)(428,251){15}
//: {16}(415,224)(400,224){17}
//: {18}(398,222)(398,212)(408,212)(408,251){19}
//: {20}(396,224)(380,224){21}
//: {22}(378,226)(378,216)(388,216)(388,251){23}
//: {24}(376,224)(360,224){25}
//: {26}(358,226)(358,216)(368,216)(368,251){27}
//: {28}(356,224)(341,224){29}
//: {30}(339,222)(339,211)(348,211)(348,251){31}
//: {32}(337,224)(320,224){33}
//: {34}(318,226)(318,216)(328,216)(328,251){35}
//: {36}(316,224)(308,224)(308,251){37}
//: {38}(318,226)(318,251){39}
//: {40}(339,226)(339,236)(338,236)(338,251){41}
//: {42}(358,226)(358,251){43}
//: {44}(378,226)(378,251){45}
//: {46}(398,226)(398,251){47}
//: {48}(417,226)(417,236)(418,236)(418,251){49}
wire w0;    //: /sn:0 {0}(618,251)(618,203){1}
wire w1;    //: /sn:0 {0}(608,251)(608,203){1}
wire w8;    //: /sn:0 {0}(578,251)(578,203){1}
wire w18;    //: /sn:0 {0}(478,251)(478,203){1}
wire w17;    //: /sn:0 {0}(488,203)(488,251){1}
wire w11;    //: /sn:0 {0}(548,251)(548,203){1}
wire w12;    //: /sn:0 {0}(538,251)(538,203){1}
wire w10;    //: /sn:0 {0}(558,203)(558,251){1}
wire w13;    //: /sn:0 {0}(528,251)(528,203){1}
wire w9;    //: /sn:0 {0}(568,251)(568,203){1}
//: enddecls

  //: joint g4 (w19) @(468, 224) /w:[ 4 6 3 8 ]
  //: joint g8 (w19) @(378, 224) /w:[ 21 22 24 44 ]
  //: OUT g3 (Sa) @(524,346) /sn:0 /w:[ 0 ]
  assign Sa = {w19, w19, w19, w19, w19, w19, w19, w19, w19, w19, w19, w19, w19, w19, w19, w19, w19, w18, w17, w16, w15, w14, w13, w12, w11, w10, w9, w8, w7, w6, w1, w0}; //: CONCAT g2  @(463,256) /sn:0 /R:3 /w:[ 1 37 39 35 41 31 43 27 45 23 47 19 49 15 0 11 5 9 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 ] /dr:1 /tp:0 /drp:1
  assign {w19, w18, w17, w16, w15, w14, w13, w12, w11, w10, w9, w8, w7, w6, w1, w0} = E; //: CONCAT g1  @(543,198) /sn:0 /R:1 /w:[ 7 1 0 1 1 1 1 1 1 0 1 1 1 1 1 1 1 ] /dr:0 /tp:0 /drp:0
  //: joint g11 (w19) @(437, 224) /w:[ 2 10 12 1 ]
  //: joint g10 (w19) @(417, 224) /w:[ 13 14 16 48 ]
  //: joint g6 (w19) @(339, 224) /w:[ 29 30 32 40 ]
  //: joint g7 (w19) @(358, 224) /w:[ 25 26 28 42 ]
  //: joint g9 (w19) @(398, 224) /w:[ 17 18 20 46 ]
  //: joint g5 (w19) @(318, 224) /w:[ 33 34 36 38 ]
  //: IN g0 (E) @(386,124) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin Mux3
module Mux3(E4, E0, C0, C1, C2, E7, E6, E2, E5, E3, E1, Sal);
//: interface  /sz:(52, 85) /bd:[ Ti0>C2(20/52) Ti1>C1(31/52) Ti2>C0(42/52) Li0>E7(78/85) Li1>E6(68/85) Li2>E5(57/85) Li3>E4(47/85) Li4>E3(38/85) Li5>E2(27/85) Li6>E1(19/85) Li7>E0(7/85) Ro0<Sal(41/85) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input E7;    //: /sn:0 {0}(502,399)(292,399)(292,410)(277,410){1}
input C0;    //: /sn:0 {0}(422,116)(422,174){1}
//: {2}(424,176)(501,176){3}
//: {4}(422,178)(422,202){5}
//: {6}(424,204)(502,204){7}
//: {8}(422,206)(422,232){9}
//: {10}(424,234)(502,234){11}
//: {12}(422,236)(422,264){13}
//: {14}(424,266)(434,266)(434,267)(502,267){15}
//: {16}(422,268)(422,300){17}
//: {18}(424,302)(434,302)(434,301)(503,301){19}
//: {20}(422,304)(422,333){21}
//: {22}(424,335)(434,335)(434,336)(503,336){23}
//: {24}(422,337)(422,367){25}
//: {26}(424,369)(434,369)(434,370)(503,370){27}
//: {28}(422,371)(422,404)(502,404){29}
input E1;    //: /sn:0 {0}(502,199)(288,199)(288,213)(273,213){1}
input E2;    //: /sn:0 {0}(502,229)(290,229)(290,248)(275,248){1}
input E0;    //: /sn:0 {0}(501,171)(287,171)(287,180)(272,180){1}
input C2;    //: /sn:0 {0}(501,186)(389,186)(389,184)(379,184){1}
//: {2}(377,182)(377,116){3}
//: {4}(377,186)(377,211){5}
//: {6}(379,213)(389,213)(389,214)(502,214){7}
//: {8}(377,215)(377,243){9}
//: {10}(379,245)(389,245)(389,244)(502,244){11}
//: {12}(377,247)(377,275){13}
//: {14}(379,277)(502,277){15}
//: {16}(377,279)(377,310){17}
//: {18}(379,312)(389,312)(389,311)(503,311){19}
//: {20}(377,314)(377,342){21}
//: {22}(379,344)(389,344)(389,346)(503,346){23}
//: {24}(377,346)(377,376){25}
//: {26}(379,378)(389,378)(389,380)(503,380){27}
//: {28}(377,380)(377,412)(389,412)(389,414)(502,414){29}
output Sal;    //: /sn:0 {0}(639,287)(731,287)(731,291)(741,291){1}
input E4;    //: /sn:0 {0}(503,296)(286,296)(286,314)(271,314){1}
input E3;    //: /sn:0 {0}(502,262)(288,262)(288,277)(273,277){1}
input E5;    //: /sn:0 {0}(503,331)(288,331)(288,349)(273,349){1}
input E6;    //: /sn:0 {0}(503,365)(291,365)(291,378)(276,378){1}
input C1;    //: /sn:0 {0}(503,375)(410,375)(410,373)(400,373){1}
//: {2}(398,371)(398,344){3}
//: {4}(400,342)(410,342)(410,341)(503,341){5}
//: {6}(398,340)(398,305){7}
//: {8}(400,303)(410,303)(410,306)(503,306){9}
//: {10}(398,301)(398,272){11}
//: {12}(400,270)(410,270)(410,272)(502,272){13}
//: {14}(398,268)(398,238){15}
//: {16}(400,236)(410,236)(410,239)(502,239){17}
//: {18}(398,234)(398,211){19}
//: {20}(400,209)(502,209){21}
//: {22}(398,207)(398,181){23}
//: {24}(400,179)(410,179)(410,181)(501,181){25}
//: {26}(398,177)(398,116){27}
//: {28}(398,375)(398,409)(502,409){29}
wire w14;    //: /sn:0 {0}(524,303)(583,303)(583,290)(618,290){1}
wire w23;    //: /sn:0 {0}(523,406)(603,406)(603,305)(618,305){1}
wire w20;    //: /sn:0 {0}(524,372)(597,372)(597,300)(618,300){1}
wire w8;    //: /sn:0 {0}(523,236)(589,236)(589,280)(618,280){1}
wire w17;    //: /sn:0 {0}(524,338)(591,338)(591,295)(618,295){1}
wire w11;    //: /sn:0 {0}(523,269)(584,269)(584,285)(618,285){1}
wire w2;    //: /sn:0 {0}(522,178)(603,178)(603,270)(618,270){1}
wire w5;    //: /sn:0 {0}(523,206)(596,206)(596,275)(618,275){1}
//: enddecls

  //: IN g8 (E4) @(269,314) /sn:0 /w:[ 1 ]
  //: IN g4 (E0) @(270,180) /sn:0 /w:[ 1 ]
  //: joint g34 (C1) @(398, 342) /w:[ 4 6 -1 3 ]
  _GGAND4 #(10) g13 (.I0(E1), .I1(C0), .I2(!C1), .I3(!C2), .Z(w5));   //: @(513,206) /sn:0 /w:[ 0 7 21 7 0 ]
  //: IN g3 (C0) @(422,114) /sn:0 /R:3 /w:[ 0 ]
  //: IN g2 (C1) @(398,114) /sn:0 /R:3 /w:[ 27 ]
  //: IN g1 (C2) @(377,114) /sn:0 /R:3 /w:[ 3 ]
  _GGAND4 #(10) g16 (.I0(E4), .I1(!C0), .I2(!C1), .I3(C2), .Z(w14));   //: @(514,303) /sn:0 /w:[ 0 19 9 19 0 ]
  //: IN g11 (E7) @(275,410) /sn:0 /w:[ 1 ]
  //: IN g10 (E6) @(274,378) /sn:0 /w:[ 1 ]
  //: joint g32 (C1) @(398, 270) /w:[ 12 14 -1 11 ]
  //: joint g27 (C0) @(422, 369) /w:[ 26 25 -1 28 ]
  _GGAND4 #(10) g19 (.I0(E7), .I1(C0), .I2(C1), .I3(C2), .Z(w23));   //: @(513,406) /sn:0 /w:[ 0 29 29 29 0 ]
  //: joint g38 (C2) @(377, 378) /w:[ 26 25 -1 28 ]
  //: IN g6 (E2) @(273,248) /sn:0 /w:[ 1 ]
  //: IN g9 (E5) @(271,349) /sn:0 /w:[ 1 ]
  //: IN g7 (E3) @(271,277) /sn:0 /w:[ 1 ]
  //: joint g31 (C1) @(398, 236) /w:[ 16 18 -1 15 ]
  _GGOR8 #(18) g20 (.I0(w2), .I1(w5), .I2(w8), .I3(w11), .I4(w14), .I5(w17), .I6(w20), .I7(w23), .Z(Sal));   //: @(629,287) /sn:0 /w:[ 1 1 1 1 1 1 1 1 0 ]
  _GGAND4 #(10) g15 (.I0(E3), .I1(C0), .I2(C1), .I3(!C2), .Z(w11));   //: @(513,269) /sn:0 /w:[ 0 15 13 15 0 ]
  //: joint g39 (C2) @(377, 344) /w:[ 22 21 -1 24 ]
  //: joint g43 (C2) @(377, 213) /w:[ 6 5 -1 8 ]
  //: joint g29 (C1) @(398, 179) /w:[ 24 26 -1 23 ]
  //: joint g25 (C0) @(422, 302) /w:[ 18 17 -1 20 ]
  _GGAND4 #(10) g17 (.I0(E5), .I1(C0), .I2(!C1), .I3(C2), .Z(w17));   //: @(514,338) /sn:0 /w:[ 0 23 5 23 0 ]
  //: joint g42 (C2) @(377, 245) /w:[ 10 9 -1 12 ]
  _GGAND4 #(10) g14 (.I0(E2), .I1(!C0), .I2(C1), .I3(!C2), .Z(w8));   //: @(513,236) /sn:0 /w:[ 0 11 17 11 0 ]
  //: IN g5 (E1) @(271,213) /sn:0 /w:[ 1 ]
  //: joint g44 (C2) @(377, 184) /w:[ 1 2 -1 4 ]
  //: joint g24 (C0) @(422, 266) /w:[ 14 13 -1 16 ]
  //: joint g21 (C0) @(422, 176) /w:[ 2 1 -1 4 ]
  //: joint g41 (C2) @(377, 277) /w:[ 14 13 -1 16 ]
  //: joint g23 (C0) @(422, 234) /w:[ 10 9 -1 12 ]
  //: joint g40 (C2) @(377, 312) /w:[ 18 17 -1 20 ]
  //: joint g35 (C1) @(398, 373) /w:[ 1 2 -1 28 ]
  //: joint g26 (C0) @(422, 335) /w:[ 22 21 -1 24 ]
  //: joint g22 (C0) @(422, 204) /w:[ 6 5 -1 8 ]
  //: OUT g0 (Sal) @(738,291) /sn:0 /w:[ 1 ]
  _GGAND4 #(10) g18 (.I0(E6), .I1(!C0), .I2(C1), .I3(C2), .Z(w20));   //: @(514,372) /sn:0 /w:[ 0 27 0 27 0 ]
  _GGAND4 #(10) g12 (.I0(E0), .I1(!C0), .I2(!C1), .I3(!C2), .Z(w2));   //: @(512,178) /sn:0 /w:[ 0 3 25 0 0 ]
  //: joint g33 (C1) @(398, 303) /w:[ 8 10 -1 7 ]
  //: joint g30 (C1) @(398, 209) /w:[ 20 22 -1 19 ]

endmodule
//: /netlistEnd

//: /netlistBegin Mux2x3
module Mux2x3(C, E1, Sa, E0, E2, E3);
//: interface  /sz:(40, 96) /bd:[ Ti0>C[1:0](19/40) Li0>E0[2:0](16/96) Li1>E1[2:0](33/96) Li2>E2[2:0](57/96) Li3>E3[2:0](78/96) Ro0<Sa[2:0](55/96) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [2:0] E1;    //: /sn:0 {0}(#:226,186)(167,186)(167,182)(#:152,182){1}
input [2:0] E2;    //: /sn:0 {0}(#:166,265)(208,265)(208,263)(#:227,263){1}
input [2:0] E0;    //: /sn:0 {0}(#:238,113)(#:149,113){1}
output [2:0] Sa;    //: /sn:0 {0}(589,251)(#:519,251){1}
input [1:0] C;    //: /sn:0 {0}(#:475,22)(511,22)(#:511,71){1}
input [2:0] E3;    //: /sn:0 {0}(#:164,345)(223,345)(223,344)(#:234,344){1}
supply0 w2;    //: /sn:0 {0}(347,403)(347,426){1}
//: {2}(349,428)(367,428)(367,403){3}
//: {4}(345,428)(328,428){5}
//: {6}(326,426)(326,416)(327,416)(327,403){7}
//: {8}(324,428)(260,428){9}
//: {10}(258,426)(258,366){11}
//: {12}(260,364)(285,364){13}
//: {14}(258,362)(258,289){15}
//: {16}(260,287)(284,287){17}
//: {18}(258,285)(258,212){19}
//: {20}(260,210)(283,210){21}
//: {22}(258,208)(258,133)(261,133){23}
//: {24}(265,133)(285,133){25}
//: {26}(263,131)(263,86)(496,86)(496,102){27}
//: {28}(263,135)(263,143)(285,143){29}
//: {30}(260,210)(250,210)(250,220)(283,220){31}
//: {32}(260,287)(250,287)(250,297)(284,297){33}
//: {34}(256,364)(246,364)(246,374)(285,374){35}
//: {36}(258,430)(258,465){37}
//: {38}(326,430)(326,440)(337,440)(337,403){39}
//: {40}(347,426)(347,436)(357,436)(357,403){41}
wire [4:0] w6;    //: /sn:0 {0}(#:375,210)(311,210)(311,277)(#:290,277){1}
wire [4:0] w7;    //: /sn:0 {0}(#:375,194)(304,194)(304,200)(#:289,200){1}
wire w14;    //: /sn:0 {0}(513,251)(464,251){1}
wire w16;    //: /sn:0 {0}(513,261)(464,261){1}
wire w15;    //: /sn:0 {0}(244,103)(285,103){1}
wire w19;    //: /sn:0 {0}(244,113)(285,113){1}
wire w38;    //: /sn:0 {0}(284,257)(248,257)(248,253)(233,253){1}
wire [2:0] w0;    //: /sn:0 {0}(#:506,108)(506,115)(396,115)(#:396,161){1}
wire w21;    //: /sn:0 {0}(285,123)(244,123){1}
wire w28;    //: /sn:0 {0}(283,180)(247,180)(247,176)(232,176){1}
wire [4:0] w1;    //: /sn:0 {0}(#:375,305)(349,305){1}
//: {2}(347,303)(347,287){3}
//: {4}(349,285)(359,285)(359,284)(#:375,284){5}
//: {6}(347,283)(347,266){7}
//: {8}(349,264)(359,264)(359,266)(#:375,266){9}
//: {10}(347,262)(347,249)(#:375,249){11}
//: {12}(347,307)(#:347,397){13}
wire [4:0] w8;    //: /sn:0 {0}(#:291,123)(360,123)(360,178)(#:375,178){1}
wire w18;    //: /sn:0 {0}(464,281)(479,281){1}
wire w40;    //: /sn:0 {0}(284,277)(248,277)(248,273)(233,273){1}
wire w30;    //: /sn:0 {0}(283,200)(247,200)(247,196)(232,196){1}
wire w17;    //: /sn:0 {0}(464,271)(479,271){1}
wire w11;    //: /sn:0 {0}(506,77)(506,102){1}
wire w12;    //: /sn:0 {0}(513,241)(464,241){1}
wire w49;    //: /sn:0 {0}(285,344)(240,344){1}
wire w10;    //: /sn:0 {0}(516,77)(516,102){1}
wire [4:0] w5;    //: /sn:0 {0}(#:375,226)(327,226)(327,354)(#:291,354){1}
wire w48;    //: /sn:0 {0}(240,334)(285,334){1}
wire w29;    //: /sn:0 {0}(283,190)(247,190)(247,186)(232,186){1}
wire [4:0] w9;    //: /sn:0 {0}(#:458,261)(#:417,261){1}
wire w50;    //: /sn:0 {0}(285,354)(240,354){1}
wire w39;    //: /sn:0 {0}(233,263)(269,263)(269,267)(284,267){1}
//: enddecls

  assign {w18, w17, w16, w14, w12} = w9; //: CONCAT g4  @(459,261) /sn:0 /R:2 /w:[ 0 0 1 1 1 0 ] /dr:0 /tp:0 /drp:0
  assign {w21, w19, w15} = E0; //: CONCAT g8  @(239,113) /sn:0 /R:2 /w:[ 1 0 0 0 ] /dr:0 /tp:0 /drp:0
  //: IN g3 (C) @(473,22) /sn:0 /w:[ 0 ]
  assign {w50, w49, w48} = E3; //: CONCAT g13  @(235,344) /sn:0 /R:2 /w:[ 1 1 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w11, w10} = C; //: CONCAT g2  @(511,72) /sn:0 /R:1 /w:[ 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign w0 = {w2, w11, w10}; //: CONCAT g1  @(506,107) /sn:0 /R:3 /w:[ 0 27 1 1 ] /dr:1 /tp:0 /drp:1
  assign {w40, w39, w38} = E2; //: CONCAT g11  @(228,263) /sn:0 /R:2 /w:[ 1 0 1 1 ] /dr:0 /tp:0 /drp:0
  //: IN g16 (E1) @(150,182) /sn:0 /w:[ 1 ]
  assign w7 = {w2, w2, w30, w29, w28}; //: CONCAT g10  @(288,200) /sn:0 /w:[ 1 31 21 0 0 0 ] /dr:1 /tp:0 /drp:1
  //: joint g28 (w2) @(258, 428) /w:[ 9 10 -1 36 ]
  assign w1 = {w2, w2, w2, w2, w2}; //: CONCAT g19  @(347,398) /sn:0 /R:1 /w:[ 13 7 39 0 41 3 ] /dr:0 /tp:0 /drp:1
  //: joint g27 (w2) @(258, 364) /w:[ 12 14 34 11 ]
  //: OUT g6 (Sa) @(586,251) /sn:0 /w:[ 0 ]
  assign w8 = {w2, w2, w21, w19, w15}; //: CONCAT g7  @(290,123) /sn:0 /w:[ 0 29 25 0 1 1 ] /dr:1 /tp:0 /drp:1
  assign {w30, w29, w28} = E1; //: CONCAT g9  @(227,186) /sn:0 /R:2 /w:[ 1 1 1 0 ] /dr:0 /tp:0 /drp:0
  //: IN g15 (E0) @(147,113) /sn:0 /w:[ 1 ]
  //: joint g20 (w1) @(347, 264) /w:[ 8 10 -1 7 ]
  //: IN g17 (E2) @(164,265) /sn:0 /w:[ 0 ]
  //: joint g25 (w2) @(258, 210) /w:[ 20 22 30 19 ]
  //: joint g29 (w2) @(326, 428) /w:[ 5 6 8 38 ]
  assign Sa = {w16, w14, w12}; //: CONCAT g5  @(518,251) /sn:0 /w:[ 1 0 0 0 ] /dr:1 /tp:0 /drp:1
  assign w5 = {w2, w2, w50, w49, w48}; //: CONCAT g14  @(290,354) /sn:0 /w:[ 1 35 13 0 0 1 ] /dr:1 /tp:0 /drp:1
  //: joint g21 (w1) @(347, 285) /w:[ 4 6 -1 3 ]
  //: joint g24 (w2) @(263, 133) /w:[ 24 26 23 28 ]
  //: GROUND g23 (w2) @(258,471) /sn:0 /w:[ 37 ]
  Mux3x5 g0 (.C(w0), .E0(w8), .E1(w7), .E2(w6), .E3(w5), .E4(w1), .E5(w1), .E6(w1), .E7(w1), .Sa(w9));   //: @(376, 162) /sz:(40, 160) /sn:0 /p:[ Ti0>1 Li0>1 Li1>0 Li2>0 Li3>0 Li4>11 Li5>9 Li6>5 Li7>0 Ro0<1 ]
  //: joint g22 (w1) @(347, 305) /w:[ 1 2 -1 12 ]
  //: joint g26 (w2) @(258, 287) /w:[ 16 18 32 15 ]
  assign w6 = {w2, w2, w40, w39, w38}; //: CONCAT g12  @(289,277) /sn:0 /w:[ 1 33 17 0 1 0 ] /dr:1 /tp:0 /drp:1
  //: IN g18 (E3) @(162,345) /sn:0 /w:[ 0 ]
  //: joint g30 (w2) @(347, 428) /w:[ 2 1 4 40 ]

endmodule
//: /netlistEnd

//: /netlistBegin Transicion
module Transicion(E0, E4, Q1, D0, E2, E3, D3, Q0, Q3, Q2, E5, D2, D1, E1);
//: interface  /sz:(90, 120) /bd:[ Ti0>Q3(19/90) Ti1>Q2(37/90) Ti2>Q1(56/90) Ti3>Q0(73/90) Li0>E5(103/120) Li1>E4(89/120) Li2>E3(76/120) Li3>E2(59/120) Li4>E1(43/120) Li5>E0(29/120) Ro0<D3(92/120) Ro1<D2(70/120) Ro2<D1(46/120) Ro3<D0(25/120) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input Q0;    //: /sn:0 {0}(323,951)(92,951){1}
//: {2}(90,949)(90,881){3}
//: {4}(92,879)(325,879){5}
//: {6}(90,877)(90,770){7}
//: {8}(92,768)(326,768){9}
//: {10}(90,766)(90,741){11}
//: {12}(92,739)(102,739)(102,738)(325,738){13}
//: {14}(90,737)(90,673){15}
//: {16}(92,671)(102,671)(102,672)(325,672){17}
//: {18}(90,669)(90,610){19}
//: {20}(92,608)(102,608)(102,610)(326,610){21}
//: {22}(90,606)(90,525){23}
//: {24}(92,523)(102,523)(102,524)(318,524){25}
//: {26}(90,521)(90,489){27}
//: {28}(92,487)(102,487)(102,488)(317,488){29}
//: {30}(90,485)(90,430){31}
//: {32}(92,428)(102,428)(102,426)(319,426){33}
//: {34}(90,426)(90,381){35}
//: {36}(92,379)(102,379)(102,380)(323,380){37}
//: {38}(90,377)(90,290){39}
//: {40}(92,288)(102,288)(102,290)(427,290){41}
//: {42}(90,286)(90,231){43}
//: {44}(92,229)(102,229)(102,231)(427,231){45}
//: {46}(90,227)(90,174){47}
//: {48}(92,172)(428,172){49}
//: {50}(90,170)(90,140){51}
//: {52}(92,138)(102,138)(102,139)(427,139){53}
//: {54}(90,136)(90,85){55}
//: {56}(92,83)(102,83)(102,84)(427,84){57}
//: {58}(90,81)(90,34){59}
//: {60}(90,953)(90,1115){61}
input E1;    //: /sn:0 {0}(214,1109)(214,926){1}
//: {2}(216,924)(226,924)(226,926)(323,926){3}
//: {4}(214,922)(214,857){5}
//: {6}(216,855)(226,855)(226,854)(325,854){7}
//: {8}(214,853)(214,715){9}
//: {10}(216,713)(325,713){11}
//: {12}(214,711)(214,649){13}
//: {14}(216,647)(325,647){15}
//: {16}(214,645)(214,592){17}
//: {18}(216,590)(326,590){19}
//: {20}(214,588)(214,468){21}
//: {22}(216,466)(226,466)(226,463)(317,463){23}
//: {24}(214,464)(214,355){25}
//: {26}(216,353)(226,353)(226,355)(323,355){27}
//: {28}(214,351)(214,268){29}
//: {30}(216,266)(301,266)(301,265)(427,265){31}
//: {32}(214,264)(214,207){33}
//: {34}(216,205)(226,205)(226,206)(427,206){35}
//: {36}(214,203)(214,117){37}
//: {38}(216,115)(226,115)(226,114)(427,114){39}
//: {40}(214,113)(214,34){41}
output D2;    //: /sn:0 {0}(452,689)(515,689)(515,690)(530,690){1}
output D1;    //: /sn:0 {0}(555,453)(446,453){1}
input E2;    //: /sn:0 {0}(323,931)(207,931)(207,930)(197,930){1}
//: {2}(195,928)(195,862){3}
//: {4}(197,860)(207,860)(207,859)(325,859){5}
//: {6}(195,858)(195,718){7}
//: {8}(197,716)(207,716)(207,718)(325,718){9}
//: {10}(195,714)(195,653){11}
//: {12}(197,651)(207,651)(207,652)(325,652){13}
//: {14}(195,649)(195,597){15}
//: {16}(197,595)(326,595){17}
//: {18}(195,593)(195,469){19}
//: {20}(197,467)(207,467)(207,468)(317,468){21}
//: {22}(195,465)(195,359){23}
//: {24}(197,357)(207,357)(207,360)(323,360){25}
//: {26}(195,355)(195,273){27}
//: {28}(197,271)(207,271)(207,270)(427,270){29}
//: {30}(195,269)(195,212){31}
//: {32}(197,210)(207,210)(207,211)(427,211){33}
//: {34}(195,208)(195,120){35}
//: {36}(197,118)(207,118)(207,119)(427,119){37}
//: {38}(195,116)(195,34){39}
//: {40}(195,932)(195,1107){41}
input E0;    //: /sn:0 {0}(427,109)(247,109)(247,108)(237,108){1}
//: {2}(235,106)(235,34){3}
//: {4}(235,110)(235,199){5}
//: {6}(237,201)(427,201){7}
//: {8}(235,203)(235,255){9}
//: {10}(237,257)(304,257)(304,260)(427,260){11}
//: {12}(235,259)(235,346){13}
//: {14}(237,348)(247,348)(247,350)(323,350){15}
//: {16}(235,350)(235,455){17}
//: {18}(237,457)(247,457)(247,458)(317,458){19}
//: {20}(235,459)(235,581){21}
//: {22}(237,583)(247,583)(247,585)(326,585){23}
//: {24}(235,585)(235,640){25}
//: {26}(237,642)(325,642){27}
//: {28}(235,644)(235,706){29}
//: {30}(237,708)(325,708){31}
//: {32}(235,710)(235,848){33}
//: {34}(237,850)(247,850)(247,849)(325,849){35}
//: {36}(235,852)(235,922){37}
//: {38}(237,924)(247,924)(247,921)(323,921){39}
//: {40}(235,926)(235,1109){41}
output D0;    //: /sn:0 {0}(578,176)(643,176)(643,175)(658,175){1}
output D3;    //: /sn:0 {0}(507,920)(447,920)(447,918)(432,918){1}
input Q1;    //: /sn:0 {0}(323,956)(76,956){1}
//: {2}(74,954)(74,884){3}
//: {4}(76,882)(86,882)(86,884)(325,884){5}
//: {6}(74,880)(74,773){7}
//: {8}(76,771)(86,771)(86,773)(326,773){9}
//: {10}(74,769)(74,744){11}
//: {12}(76,742)(86,742)(86,743)(325,743){13}
//: {14}(74,740)(74,679){15}
//: {16}(76,677)(325,677){17}
//: {18}(74,675)(74,617){19}
//: {20}(76,615)(326,615){21}
//: {22}(74,613)(74,528){23}
//: {24}(76,526)(86,526)(86,529)(318,529){25}
//: {26}(74,524)(74,493){27}
//: {28}(76,491)(86,491)(86,493)(317,493){29}
//: {30}(74,489)(74,434){31}
//: {32}(76,432)(86,432)(86,431)(319,431){33}
//: {34}(74,430)(74,386){35}
//: {36}(76,384)(86,384)(86,385)(323,385){37}
//: {38}(74,382)(74,298){39}
//: {40}(76,296)(86,296)(86,295)(427,295){41}
//: {42}(74,294)(74,238){43}
//: {44}(76,236)(427,236){45}
//: {46}(74,234)(74,179){47}
//: {48}(76,177)(428,177){49}
//: {50}(74,175)(74,145){51}
//: {52}(76,143)(86,143)(86,144)(427,144){53}
//: {54}(74,141)(74,90){55}
//: {56}(76,88)(86,88)(86,89)(427,89){57}
//: {58}(74,86)(74,34){59}
//: {60}(74,958)(74,1116){61}
input E4;    //: /sn:0 {0}(323,941)(166,941)(166,940)(156,940){1}
//: {2}(154,938)(154,869){3}
//: {4}(156,867)(166,867)(166,869)(325,869){5}
//: {6}(154,865)(154,727){7}
//: {8}(156,725)(166,725)(166,728)(325,728){9}
//: {10}(154,723)(154,665){11}
//: {12}(156,663)(166,663)(166,662)(325,662){13}
//: {14}(154,661)(154,600){15}
//: {16}(156,598)(166,598)(166,600)(326,600){17}
//: {18}(154,596)(154,478){19}
//: {20}(156,476)(166,476)(166,478)(317,478){21}
//: {22}(154,474)(154,369){23}
//: {24}(156,367)(166,367)(166,370)(323,370){25}
//: {26}(154,365)(154,281){27}
//: {28}(156,279)(166,279)(166,280)(427,280){29}
//: {30}(154,277)(154,222){31}
//: {32}(156,220)(166,220)(166,221)(427,221){33}
//: {34}(154,218)(154,130){35}
//: {36}(156,128)(166,128)(166,129)(427,129){37}
//: {38}(154,126)(154,34){39}
//: {40}(154,942)(154,1105){41}
input Q3;    //: /sn:0 {0}(323,966)(49,966)(49,967)(39,967){1}
//: {2}(37,965)(37,894){3}
//: {4}(39,892)(49,892)(49,894)(325,894){5}
//: {6}(37,890)(37,784){7}
//: {8}(39,782)(49,782)(49,783)(326,783){9}
//: {10}(37,780)(37,753){11}
//: {12}(39,751)(49,751)(49,753)(325,753){13}
//: {14}(37,749)(37,689){15}
//: {16}(39,687)(325,687){17}
//: {18}(37,685)(37,628){19}
//: {20}(39,626)(49,626)(49,625)(326,625){21}
//: {22}(37,624)(37,537){23}
//: {24}(39,535)(49,535)(49,539)(318,539){25}
//: {26}(37,533)(37,504){27}
//: {28}(39,502)(49,502)(49,503)(317,503){29}
//: {30}(37,500)(37,443){31}
//: {32}(39,441)(319,441){33}
//: {34}(37,439)(37,395){35}
//: {36}(39,393)(49,393)(49,395)(323,395){37}
//: {38}(37,391)(37,305){39}
//: {40}(39,303)(49,303)(49,305)(427,305){41}
//: {42}(37,301)(37,246){43}
//: {44}(39,244)(49,244)(49,246)(427,246){45}
//: {46}(37,242)(37,189){47}
//: {48}(39,187)(428,187){49}
//: {50}(37,185)(37,154){51}
//: {52}(39,152)(49,152)(49,154)(427,154){53}
//: {54}(37,150)(37,103){55}
//: {56}(39,101)(49,101)(49,99)(427,99){57}
//: {58}(37,99)(37,34){59}
//: {60}(37,969)(37,1115){61}
input E3;    //: /sn:0 {0}(323,936)(187,936)(187,933)(177,933){1}
//: {2}(175,931)(175,866){3}
//: {4}(177,864)(325,864){5}
//: {6}(175,862)(175,724){7}
//: {8}(177,722)(187,722)(187,723)(325,723){9}
//: {10}(175,720)(175,659){11}
//: {12}(177,657)(325,657){13}
//: {14}(175,655)(175,477){15}
//: {16}(177,475)(187,475)(187,473)(317,473){17}
//: {18}(175,473)(175,366){19}
//: {20}(177,364)(187,364)(187,365)(323,365){21}
//: {22}(175,362)(175,276){23}
//: {24}(177,274)(187,274)(187,275)(427,275){25}
//: {26}(175,272)(175,219){27}
//: {28}(177,217)(187,217)(187,216)(427,216){29}
//: {30}(175,215)(175,126){31}
//: {32}(177,124)(427,124){33}
//: {34}(175,122)(175,34){35}
//: {36}(175,935)(175,1109){37}
input E5;    //: /sn:0 {0}(323,946)(144,946)(144,943)(134,943){1}
//: {2}(132,941)(132,874){3}
//: {4}(134,872)(144,872)(144,874)(325,874){5}
//: {6}(132,870)(132,734){7}
//: {8}(134,732)(144,732)(144,733)(325,733){9}
//: {10}(132,730)(132,668){11}
//: {12}(134,666)(144,666)(144,667)(325,667){13}
//: {14}(132,664)(132,608){15}
//: {16}(134,606)(144,606)(144,605)(326,605){17}
//: {18}(132,604)(132,484){19}
//: {20}(134,482)(144,482)(144,483)(317,483){21}
//: {22}(132,480)(132,377){23}
//: {24}(134,375)(323,375){25}
//: {26}(132,373)(132,285){27}
//: {28}(134,283)(144,283)(144,285)(427,285){29}
//: {30}(132,281)(132,226){31}
//: {32}(134,224)(144,224)(144,226)(427,226){33}
//: {34}(132,222)(132,134){35}
//: {36}(134,132)(144,132)(144,134)(427,134){37}
//: {38}(132,130)(132,34){39}
//: {40}(132,945)(132,1107){41}
input Q2;    //: /sn:0 {0}(323,961)(66,961)(66,960)(56,960){1}
//: {2}(54,958)(54,889){3}
//: {4}(56,887)(66,887)(66,889)(325,889){5}
//: {6}(54,885)(54,779){7}
//: {8}(56,777)(66,777)(66,778)(326,778){9}
//: {10}(54,775)(54,748){11}
//: {12}(56,746)(66,746)(66,748)(325,748){13}
//: {14}(54,744)(54,683){15}
//: {16}(56,681)(66,681)(66,682)(325,682){17}
//: {18}(54,679)(54,622){19}
//: {20}(56,620)(326,620){21}
//: {22}(54,618)(54,532){23}
//: {24}(56,530)(66,530)(66,534)(318,534){25}
//: {26}(54,528)(54,499){27}
//: {28}(56,497)(66,497)(66,498)(317,498){29}
//: {30}(54,495)(54,437){31}
//: {32}(56,435)(66,435)(66,436)(319,436){33}
//: {34}(54,433)(54,393){35}
//: {36}(56,391)(66,391)(66,390)(323,390){37}
//: {38}(54,389)(54,302){39}
//: {40}(56,300)(427,300){41}
//: {42}(54,298)(54,242){43}
//: {44}(56,240)(66,240)(66,241)(427,241){45}
//: {46}(54,238)(54,187){47}
//: {48}(56,185)(66,185)(66,182)(428,182){49}
//: {50}(54,183)(54,151){51}
//: {52}(56,149)(427,149){53}
//: {54}(54,147)(54,98){55}
//: {56}(56,96)(66,96)(66,94)(427,94){57}
//: {58}(54,94)(54,34){59}
//: {60}(54,962)(54,1115){61}
wire w6;    //: /sn:0 {0}(557,176)(464,176)(464,179)(449,179){1}
wire w7;    //: /sn:0 {0}(425,456)(353,456)(353,480)(338,480){1}
wire w14;    //: /sn:0 {0}(347,775)(416,775)(416,697)(431,697){1}
wire w4;    //: /sn:0 {0}(425,446)(410,446)(410,372)(344,372){1}
wire w3;    //: /sn:0 {0}(557,171)(532,171)(532,131)(448,131){1}
wire w21;    //: /sn:0 {0}(346,871)(389,871)(389,915)(411,915){1}
wire w18;    //: /sn:0 {0}(411,920)(387,920)(387,943)(344,943){1}
wire w8;    //: /sn:0 {0}(339,531)(410,531)(410,461)(425,461){1}
wire w11;    //: /sn:0 {0}(431,687)(361,687)(361,664)(346,664){1}
wire w12;    //: /sn:0 {0}(448,282)(542,282)(542,186)(557,186){1}
wire w2;    //: /sn:0 {0}(448,91)(542,91)(542,166)(557,166){1}
wire w10;    //: /sn:0 {0}(347,605)(416,605)(416,682)(431,682){1}
wire w13;    //: /sn:0 {0}(431,692)(361,692)(361,730)(346,730){1}
wire w5;    //: /sn:0 {0}(425,451)(355,451)(355,433)(340,433){1}
wire w9;    //: /sn:0 {0}(557,181)(476,181)(476,223)(448,223){1}
//: enddecls

  //: IN g4 (E0) @(235,32) /sn:0 /R:3 /w:[ 3 ]
  //: IN g8 (E4) @(154,32) /sn:0 /R:3 /w:[ 39 ]
  //: joint g140 (E0) @(235, 924) /w:[ 38 37 -1 40 ]
  //: joint g13 (Q2) @(54, 96) /w:[ 56 58 -1 55 ]
  //: joint g37 (E4) @(154, 220) /w:[ 32 34 -1 31 ]
  _GGAND10 #(22) g55 (.I0(!E0), .I1(!E1), .I2(!E2), .I3(!E3), .I4(!E4), .I5(!E5), .I6(Q0), .I7(!Q1), .I8(!Q2), .I9(!Q3), .Z(w4));   //: @(334,372) /sn:0 /w:[ 15 27 25 21 25 25 37 37 37 37 1 ]
  //: joint g58 (E2) @(195, 357) /w:[ 24 26 -1 23 ]
  //: joint g139 (Q3) @(37, 892) /w:[ 4 6 -1 3 ]
  //: joint g112 (E1) @(214, 713) /w:[ 10 12 -1 9 ]
  //: joint g76 (E3) @(175, 475) /w:[ 16 18 -1 15 ]
  //: joint g111 (E0) @(235, 708) /w:[ 30 29 -1 32 ]
  //: IN g1 (Q1) @(74,32) /sn:0 /R:3 /w:[ 59 ]
  //: joint g64 (Q2) @(54, 391) /w:[ 36 38 -1 35 ]
  //: joint g11 (Q0) @(90, 83) /w:[ 56 58 -1 55 ]
  //: joint g130 (E0) @(235, 850) /w:[ 34 33 -1 36 ]
  _GGAND4 #(10) g121 (.I0(Q0), .I1(!Q1), .I2(Q2), .I3(!Q3), .Z(w14));   //: @(337,775) /sn:0 /w:[ 9 9 9 9 0 ]
  //: joint g28 (Q3) @(37, 152) /w:[ 52 54 -1 51 ]
  //: OUT g50 (D0) @(655,175) /sn:0 /w:[ 1 ]
  //: joint g132 (E2) @(195, 860) /w:[ 4 6 -1 3 ]
  //: joint g19 (E0) @(235, 108) /w:[ 1 2 -1 4 ]
  //: joint g113 (E2) @(195, 716) /w:[ 8 10 -1 7 ]
  _GGOR2 #(6) g150 (.I0(w21), .I1(w18), .Z(D3));   //: @(422,918) /sn:0 /w:[ 1 0 1 ]
  //: joint g146 (Q0) @(90, 951) /w:[ 1 2 -1 60 ]
  //: IN g6 (E2) @(195,32) /sn:0 /R:3 /w:[ 39 ]
  //: joint g38 (E5) @(132, 224) /w:[ 32 34 -1 31 ]
  //: joint g115 (E4) @(154, 725) /w:[ 8 10 -1 7 ]
  //: IN g7 (E3) @(175,32) /sn:0 /R:3 /w:[ 35 ]
  //: joint g53 (Q2) @(54, 300) /w:[ 40 42 -1 39 ]
  //: joint g75 (E4) @(154, 476) /w:[ 20 22 -1 19 ]
  //: joint g135 (E5) @(132, 872) /w:[ 4 6 -1 3 ]
  //: joint g20 (E1) @(214, 115) /w:[ 38 40 -1 37 ]
  //: joint g31 (Q2) @(54, 185) /w:[ 48 50 -1 47 ]
  //: joint g149 (Q3) @(37, 967) /w:[ 1 2 -1 60 ]
  //: joint g124 (Q1) @(74, 771) /w:[ 8 10 -1 7 ]
  //: joint g39 (Q0) @(90, 229) /w:[ 44 46 -1 43 ]
  //: joint g68 (Q1) @(74, 432) /w:[ 32 34 -1 31 ]
  //: joint g48 (E5) @(132, 283) /w:[ 28 30 -1 27 ]
  _GGAND10 #(22) g17 (.I0(E0), .I1(E1), .I2(!E2), .I3(!E3), .I4(!E4), .I5(E5), .I6(!Q0), .I7(!Q1), .I8(Q2), .I9(!Q3), .Z(w9));   //: @(438,223) /sn:0 /w:[ 7 35 33 29 33 33 45 45 45 45 1 ]
  //: joint g25 (Q0) @(90, 138) /w:[ 52 54 -1 51 ]
  //: joint g29 (Q0) @(90, 172) /w:[ 48 50 -1 47 ]
  //: joint g52 (Q1) @(74, 296) /w:[ 40 42 -1 39 ]
  //: joint g106 (Q0) @(90, 671) /w:[ 16 18 -1 15 ]
  //: joint g107 (Q1) @(74, 677) /w:[ 16 18 -1 15 ]
  //: joint g83 (Q0) @(90, 523) /w:[ 24 26 -1 23 ]
  //: joint g100 (E0) @(235, 642) /w:[ 26 25 -1 28 ]
  //: joint g14 (Q3) @(37, 101) /w:[ 56 58 -1 55 ]
  //: joint g44 (E1) @(214, 266) /w:[ 30 32 -1 29 ]
  //: joint g47 (E4) @(154, 279) /w:[ 28 30 -1 27 ]
  //: joint g80 (Q2) @(54, 497) /w:[ 28 30 -1 27 ]
  //: joint g94 (E5) @(132, 606) /w:[ 16 18 -1 15 ]
  //: joint g21 (E2) @(195, 118) /w:[ 36 38 -1 35 ]
  //: joint g84 (Q1) @(74, 526) /w:[ 24 26 -1 23 ]
  //: joint g105 (E5) @(132, 666) /w:[ 12 14 -1 11 ]
  //: joint g141 (E1) @(214, 924) /w:[ 2 4 -1 1 ]
  //: joint g23 (E4) @(154, 128) /w:[ 36 38 -1 35 ]
  //: joint g41 (Q2) @(54, 240) /w:[ 44 46 -1 43 ]
  //: OUT g151 (D3) @(504,920) /sn:0 /w:[ 0 ]
  //: joint g40 (Q1) @(74, 236) /w:[ 44 46 -1 43 ]
  //: joint g54 (Q3) @(37, 303) /w:[ 40 42 -1 39 ]
  //: joint g93 (E4) @(154, 598) /w:[ 16 18 -1 15 ]
  //: joint g116 (E5) @(132, 732) /w:[ 8 10 -1 7 ]
  //: joint g123 (Q2) @(54, 777) /w:[ 8 10 -1 7 ]
  //: IN g0 (Q0) @(90,32) /sn:0 /R:3 /w:[ 59 ]
  //: joint g26 (Q1) @(74, 143) /w:[ 52 54 -1 51 ]
  //: joint g46 (E3) @(175, 274) /w:[ 24 26 -1 23 ]
  //: joint g90 (E0) @(235, 583) /w:[ 22 21 -1 24 ]
  _GGAND4 #(10) g82 (.I0(Q0), .I1(!Q1), .I2(Q2), .I3(!Q3), .Z(w8));   //: @(329,531) /sn:0 /w:[ 25 25 25 25 0 ]
  //: joint g136 (E4) @(154, 867) /w:[ 4 6 -1 3 ]
  _GGAND10 #(22) g128 (.I0(!E0), .I1(!E1), .I2(E2), .I3(!E3), .I4(!E4), .I5(!E5), .I6(Q0), .I7(!Q1), .I8(!Q2), .I9(!Q3), .Z(w21));   //: @(336,871) /sn:0 /w:[ 35 7 5 5 5 5 5 5 5 5 0 ]
  //: joint g33 (E0) @(235, 201) /w:[ 6 5 -1 8 ]
  //: joint g91 (E1) @(214, 590) /w:[ 18 20 -1 17 ]
  _GGOR5 #(12) g49 (.I0(w2), .I1(w3), .I2(w6), .I3(w9), .I4(w12), .Z(D0));   //: @(568,176) /sn:0 /w:[ 1 0 0 0 1 0 ]
  //: joint g137 (Q1) @(74, 882) /w:[ 4 6 -1 3 ]
  //: joint g61 (E5) @(132, 375) /w:[ 24 26 -1 23 ]
  //: IN g3 (Q3) @(37,32) /sn:0 /R:3 /w:[ 59 ]
  //: joint g34 (E1) @(214, 205) /w:[ 34 36 -1 33 ]
  //: joint g51 (Q0) @(90, 288) /w:[ 40 42 -1 39 ]
  //: joint g86 (Q3) @(37, 535) /w:[ 24 26 -1 23 ]
  _GGAND9 #(20) g89 (.I0(E0), .I1(E1), .I2(!E2), .I3(!E4), .I4(E5), .I5(Q0), .I6(!Q1), .I7(!Q2), .I8(!Q3), .Z(w10));   //: @(337,605) /sn:0 /w:[ 23 19 17 17 17 21 21 21 21 0 ]
  //: IN g2 (Q2) @(54,32) /sn:0 /R:3 /w:[ 59 ]
  //: joint g65 (Q3) @(37, 393) /w:[ 36 38 -1 35 ]
  //: joint g77 (E5) @(132, 482) /w:[ 20 22 -1 19 ]
  _GGAND10 #(22) g110 (.I0(E0), .I1(E1), .I2(!E2), .I3(E3), .I4(!E4), .I5(E5), .I6(!Q0), .I7(!Q1), .I8(Q2), .I9(!Q3), .Z(w13));   //: @(336,730) /sn:0 /w:[ 31 11 9 9 9 9 13 13 13 13 1 ]
  //: joint g148 (Q2) @(54, 960) /w:[ 1 2 -1 60 ]
  //: joint g147 (Q1) @(74, 956) /w:[ 1 2 -1 60 ]
  //: joint g59 (E3) @(175, 364) /w:[ 20 22 -1 19 ]
  //: joint g72 (E0) @(235, 457) /w:[ 18 17 -1 20 ]
  //: joint g98 (Q3) @(37, 626) /w:[ 20 22 -1 19 ]
  _GGAND10 #(22) g99 (.I0(E0), .I1(E1), .I2(!E2), .I3(!E3), .I4(!E4), .I5(E5), .I6(!Q0), .I7(!Q1), .I8(Q2), .I9(!Q3), .Z(w11));   //: @(336,664) /sn:0 /w:[ 27 15 13 13 13 13 17 17 17 17 1 ]
  _GGAND4 #(10) g16 (.I0(!Q0), .I1(Q1), .I2(!Q2), .I3(!Q3), .Z(w6));   //: @(439,179) /sn:0 /w:[ 49 49 49 49 1 ]
  //: joint g96 (Q1) @(74, 615) /w:[ 20 22 -1 19 ]
  //: joint g103 (E3) @(175, 657) /w:[ 12 14 -1 11 ]
  //: joint g122 (Q0) @(90, 768) /w:[ 8 10 -1 7 ]
  _GGAND4 #(8) g10 (.I0(!Q0), .I1(!Q1), .I2(!Q2), .I3(!Q3), .Z(w2));   //: @(438,91) /sn:0 /w:[ 57 57 57 57 0 ]
  //: joint g78 (Q0) @(90, 487) /w:[ 28 30 -1 27 ]
  _GGOR4 #(10) g87 (.I0(w4), .I1(w5), .I2(w7), .I3(w8), .Z(D1));   //: @(436,453) /sn:0 /w:[ 0 0 0 1 1 ]
  _GGAND10 #(22) g129 (.I0(!E0), .I1(E1), .I2(!E2), .I3(!E3), .I4(!E4), .I5(!E5), .I6(Q0), .I7(!Q1), .I8(!Q2), .I9(!Q3), .Z(w18));   //: @(334,943) /sn:0 /w:[ 39 3 0 0 0 0 0 0 0 0 1 ]
  //: joint g27 (Q2) @(54, 149) /w:[ 52 54 -1 51 ]
  //: joint g32 (Q3) @(37, 187) /w:[ 48 50 -1 47 ]
  //: joint g102 (E2) @(195, 651) /w:[ 12 14 -1 11 ]
  //: joint g143 (E3) @(175, 933) /w:[ 1 2 -1 36 ]
  //: joint g69 (Q2) @(54, 435) /w:[ 32 34 -1 31 ]
  //: IN g9 (E5) @(132,32) /sn:0 /R:3 /w:[ 39 ]
  //: joint g57 (E1) @(214, 353) /w:[ 26 28 -1 25 ]
  //: joint g119 (Q2) @(54, 746) /w:[ 12 14 -1 11 ]
  //: joint g142 (E2) @(195, 930) /w:[ 1 2 -1 40 ]
  _GGAND10 #(22) g15 (.I0(!E0), .I1(E1), .I2(!E2), .I3(!E3), .I4(!E4), .I5(!E5), .I6(Q0), .I7(!Q1), .I8(!Q2), .I9(!Q3), .Z(w3));   //: @(438,131) /sn:0 /w:[ 0 39 37 33 37 37 53 53 53 53 1 ]
  _GGAND10 #(22) g71 (.I0(E0), .I1(E1), .I2(!E2), .I3(E3), .I4(!E4), .I5(E5), .I6(!Q0), .I7(!Q1), .I8(Q2), .I9(!Q3), .Z(w7));   //: @(328,480) /sn:0 /w:[ 19 23 21 17 21 21 29 29 29 29 1 ]
  //: joint g131 (E1) @(214, 855) /w:[ 6 8 -1 5 ]
  //: joint g67 (Q0) @(90, 428) /w:[ 32 34 -1 31 ]
  //: OUT g127 (D2) @(527,690) /sn:0 /w:[ 1 ]
  //: joint g43 (E0) @(235, 257) /w:[ 10 9 -1 12 ]
  //: joint g145 (E5) @(132, 943) /w:[ 1 2 -1 40 ]
  //: joint g62 (Q0) @(90, 379) /w:[ 36 38 -1 35 ]
  //: joint g73 (E1) @(214, 466) /w:[ 22 24 -1 21 ]
  //: OUT g88 (D1) @(552,453) /sn:0 /w:[ 0 ]
  //: joint g104 (E4) @(154, 663) /w:[ 12 14 -1 11 ]
  //: joint g138 (Q2) @(54, 887) /w:[ 4 6 -1 3 ]
  //: joint g42 (Q3) @(37, 244) /w:[ 44 46 -1 43 ]
  //: joint g63 (Q1) @(74, 384) /w:[ 36 38 -1 35 ]
  //: joint g74 (E2) @(195, 467) /w:[ 20 22 -1 19 ]
  //: joint g109 (Q3) @(37, 687) /w:[ 16 18 -1 15 ]
  //: joint g133 (E3) @(175, 864) /w:[ 4 6 -1 3 ]
  //: IN g5 (E1) @(214,32) /sn:0 /R:3 /w:[ 41 ]
  //: joint g56 (E0) @(235, 348) /w:[ 14 13 -1 16 ]
  //: joint g79 (Q1) @(74, 491) /w:[ 28 30 -1 27 ]
  //: joint g95 (Q0) @(90, 608) /w:[ 20 22 -1 19 ]
  //: joint g117 (Q0) @(90, 739) /w:[ 12 14 -1 11 ]
  //: joint g24 (E5) @(132, 132) /w:[ 36 38 -1 35 ]
  //: joint g36 (E3) @(175, 217) /w:[ 28 30 -1 27 ]
  //: joint g85 (Q2) @(54, 530) /w:[ 24 26 -1 23 ]
  //: joint g92 (E2) @(195, 595) /w:[ 16 18 -1 15 ]
  //: joint g144 (E4) @(154, 940) /w:[ 1 2 -1 40 ]
  //: joint g125 (Q3) @(37, 782) /w:[ 8 10 -1 7 ]
  //: joint g60 (E4) @(154, 367) /w:[ 24 26 -1 23 ]
  //: joint g81 (Q3) @(37, 502) /w:[ 28 30 -1 27 ]
  //: joint g101 (E1) @(214, 647) /w:[ 14 16 -1 13 ]
  //: joint g22 (E3) @(175, 124) /w:[ 32 34 -1 31 ]
  //: joint g35 (E2) @(195, 210) /w:[ 32 34 -1 31 ]
  //: joint g45 (E2) @(195, 271) /w:[ 28 30 -1 27 ]
  //: joint g70 (Q3) @(37, 441) /w:[ 32 34 -1 31 ]
  _GGOR4 #(10) g126 (.I0(w10), .I1(w11), .I2(w13), .I3(w14), .Z(D2));   //: @(442,689) /sn:0 /w:[ 1 0 0 1 0 ]
  _GGAND4 #(10) g66 (.I0(!Q0), .I1(Q1), .I2(!Q2), .I3(!Q3), .Z(w5));   //: @(330,433) /sn:0 /w:[ 33 33 33 33 1 ]
  //: joint g97 (Q2) @(54, 620) /w:[ 20 22 -1 19 ]
  //: joint g114 (E3) @(175, 722) /w:[ 8 10 -1 7 ]
  //: joint g120 (Q3) @(37, 751) /w:[ 12 14 -1 11 ]
  _GGAND10 #(22) g18 (.I0(E0), .I1(E1), .I2(!E2), .I3(E3), .I4(!E4), .I5(E5), .I6(!Q0), .I7(!Q1), .I8(Q2), .I9(!Q3), .Z(w12));   //: @(438,282) /sn:0 /w:[ 11 31 29 25 29 29 41 41 41 41 0 ]
  //: joint g12 (Q1) @(74, 88) /w:[ 56 58 -1 55 ]
  //: joint g30 (Q1) @(74, 177) /w:[ 48 50 -1 47 ]
  //: joint g108 (Q2) @(54, 681) /w:[ 16 18 -1 15 ]
  //: joint g134 (Q0) @(90, 879) /w:[ 4 6 -1 3 ]
  //: joint g118 (Q1) @(74, 742) /w:[ 12 14 -1 11 ]

endmodule
//: /netlistEnd

//: /netlistBegin Overflow
module Overflow(Sa, SiSa, B31, A31, R);
//: interface  /sz:(111, 43) /bd:[ Ti0>A31(42/111) Ti1>B31(63/111) Ti2>R(20/111) Ti3>SiSa(85/111) Bo0<Sa(54/111) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input A31;    //: /sn:0 {0}(286,245)(286,113){1}
//: {2}(288,111)(334,111){3}
//: {4}(338,111)(383,111){5}
//: {6}(387,111)(427,111)(427,244){7}
//: {8}(385,113)(385,245){9}
//: {10}(336,113)(336,123)(337,123)(337,246){11}
//: {12}(284,111)(130,111){13}
input SiSa;    //: /sn:0 {0}(126,190)(294,190){1}
//: {2}(298,190)(345,190){3}
//: {4}(349,190)(393,190){5}
//: {6}(397,190)(437,190)(437,244){7}
//: {8}(395,192)(395,245){9}
//: {10}(347,192)(347,246){11}
//: {12}(296,192)(296,245){13}
input R;    //: /sn:0 {0}(281,245)(281,88)(280,88)(280,78){1}
//: {2}(282,76)(327,76){3}
//: {4}(331,76)(378,76){5}
//: {6}(382,76)(422,76)(422,244){7}
//: {8}(380,78)(380,245){9}
//: {10}(329,78)(329,88)(332,88)(332,246){11}
//: {12}(278,76)(127,76){13}
output Sa;    //: /sn:0 {0}(616,416)(364,416)(364,353){1}
input B31;    //: /sn:0 {0}(126,152)(251,152)(251,151)(290,151){1}
//: {2}(294,151)(339,151){3}
//: {4}(343,151)(387,151){5}
//: {6}(391,151)(432,151)(432,244){7}
//: {8}(389,153)(389,163)(390,163)(390,245){9}
//: {10}(341,153)(341,163)(342,163)(342,246){11}
//: {12}(292,153)(292,163)(291,163)(291,245){13}
wire w11;    //: /sn:0 {0}(430,265)(430,317)(371,317)(371,332){1}
wire w12;    //: /sn:0 {0}(289,266)(289,317)(356,317)(356,332){1}
wire w2;    //: /sn:0 {0}(361,332)(361,277)(340,277)(340,267){1}
wire w5;    //: /sn:0 {0}(366,332)(366,276)(388,276)(388,266){1}
//: enddecls

  //: OUT g4 (Sa) @(613,416) /sn:0 /w:[ 0 ]
  _GGAND4 #(10) g8 (.I0(!SiSa), .I1(!B31), .I2(A31), .I3(R), .Z(w11));   //: @(430,255) /sn:0 /R:3 /w:[ 7 7 7 7 0 ]
  //: IN g3 (SiSa) @(124,190) /sn:0 /w:[ 0 ]
  //: joint g13 (R) @(380, 76) /w:[ 6 -1 5 8 ]
  //: IN g2 (B31) @(124,152) /sn:0 /w:[ 0 ]
  //: IN g1 (A31) @(128,111) /sn:0 /w:[ 13 ]
  //: joint g11 (B31) @(389, 151) /w:[ 6 -1 5 8 ]
  //: joint g16 (A31) @(336, 111) /w:[ 4 -1 3 10 ]
  //: joint g10 (SiSa) @(395, 190) /w:[ 6 -1 5 8 ]
  //: joint g19 (B31) @(292, 151) /w:[ 2 -1 1 12 ]
  _GGAND4 #(10) g6 (.I0(!SiSa), .I1(B31), .I2(A31), .I3(!R), .Z(w2));   //: @(340,257) /sn:0 /R:3 /w:[ 11 11 11 11 1 ]
  _GGAND4 #(10) g7 (.I0(SiSa), .I1(B31), .I2(!A31), .I3(R), .Z(w5));   //: @(388,256) /sn:0 /R:3 /w:[ 9 9 9 9 1 ]
  _GGOR4 #(10) g9 (.I0(w11), .I1(w5), .I2(w2), .I3(w12), .Z(Sa));   //: @(364,343) /sn:0 /R:3 /w:[ 1 0 0 1 1 ]
  //: joint g15 (B31) @(341, 151) /w:[ 4 -1 3 10 ]
  //: joint g20 (A31) @(286, 111) /w:[ 2 -1 12 1 ]
  //: joint g17 (R) @(329, 76) /w:[ 4 -1 3 10 ]
  _GGAND4 #(10) g5 (.I0(SiSa), .I1(!B31), .I2(!A31), .I3(!R), .Z(w12));   //: @(289,256) /sn:0 /R:3 /w:[ 13 13 0 0 0 ]
  //: joint g14 (SiSa) @(347, 190) /w:[ 4 -1 3 10 ]
  //: joint g21 (R) @(280, 76) /w:[ 2 -1 12 1 ]
  //: IN g0 (R) @(125,76) /sn:0 /w:[ 13 ]
  //: joint g12 (A31) @(385, 111) /w:[ 6 -1 5 8 ]
  //: joint g18 (SiSa) @(296, 190) /w:[ 2 -1 1 12 ]

endmodule
//: /netlistEnd

//: /netlistBegin n4
module n4(Sa);
//: interface  /sz:(40, 40) /bd:[ Ro0<Sa[31:0](20/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
supply0 w3;    //: /sn:0 {0}(347,113)(308,113){1}
//: {2}(306,111)(306,83)(347,83){3}
//: {4}(304,113)(291,113){5}
//: {6}(289,111)(289,73)(320,73){7}
//: {8}(324,73)(347,73){9}
//: {10}(322,75)(322,103)(347,103){11}
//: {12}(287,113)(277,113)(277,123)(347,123){13}
//: {14}(289,115)(289,141){15}
//: {16}(291,143)(347,143){17}
//: {18}(291,143)(281,143)(281,133)(347,133){19}
//: {20}(289,145)(289,161){21}
//: {22}(291,163)(347,163){23}
//: {24}(291,163)(281,163)(281,153)(347,153){25}
//: {26}(289,165)(289,181){27}
//: {28}(291,183)(347,183){29}
//: {30}(291,183)(281,183)(281,173)(347,173){31}
//: {32}(289,185)(289,200){33}
//: {34}(291,202)(301,202)(301,203)(347,203){35}
//: {36}(287,202)(277,202)(277,193)(347,193){37}
//: {38}(289,204)(289,222){39}
//: {40}(291,224)(301,224)(301,223)(347,223){41}
//: {42}(291,224)(281,224)(281,213)(347,213){43}
//: {44}(289,226)(289,242){45}
//: {46}(291,244)(301,244)(301,243)(347,243){47}
//: {48}(291,244)(281,244)(281,233)(347,233){49}
//: {50}(289,246)(289,261){51}
//: {52}(291,263)(347,263){53}
//: {54}(291,263)(281,263)(281,253)(347,253){55}
//: {56}(289,265)(289,281){57}
//: {58}(291,283)(347,283){59}
//: {60}(291,283)(281,283)(281,273)(347,273){61}
//: {62}(289,285)(289,300){63}
//: {64}(291,302)(301,302)(301,303)(347,303){65}
//: {66}(291,302)(281,302)(281,293)(347,293){67}
//: {68}(289,304)(289,320){69}
//: {70}(291,322)(301,322)(301,323)(347,323){71}
//: {72}(287,322)(277,322)(277,313)(347,313){73}
//: {74}(289,324)(289,341){75}
//: {76}(291,343)(347,343){77}
//: {78}(287,343)(277,343)(277,333)(347,333){79}
//: {80}(289,345)(289,361){81}
//: {82}(291,363)(347,363){83}
//: {84}(287,363)(277,363)(277,353)(347,353){85}
//: {86}(289,365)(289,380){87}
//: {88}(291,382)(301,382)(301,383)(347,383){89}
//: {90}(287,382)(277,382)(277,373)(347,373){91}
//: {92}(289,384)(289,432){93}
output [31:0] Sa;    //: /sn:0 {0}(394,228)(#:353,228){1}
supply1 w2;    //: /sn:0 {0}(140,47)(140,93)(347,93){1}
//: enddecls

  //: joint g8 (w3) @(289, 302) /w:[ 64 63 66 68 ]
  //: joint g4 (w3) @(289, 382) /w:[ 88 87 90 92 ]
  //: joint g13 (w3) @(289, 202) /w:[ 34 33 36 38 ]
  //: GROUND g3 (w3) @(289,438) /sn:0 /w:[ 93 ]
  //: VDD g2 (w2) @(151,47) /sn:0 /w:[ 0 ]
  //: OUT g1 (Sa) @(391,228) /sn:0 /w:[ 0 ]
  //: joint g16 (w3) @(289, 143) /w:[ 16 15 18 20 ]
  //: joint g11 (w3) @(289, 244) /w:[ 46 45 48 50 ]
  //: joint g10 (w3) @(289, 263) /w:[ 52 51 54 56 ]
  //: joint g19 (w3) @(306, 113) /w:[ 1 2 4 -1 ]
  //: joint g6 (w3) @(289, 343) /w:[ 76 75 78 80 ]
  //: joint g9 (w3) @(289, 283) /w:[ 58 57 60 62 ]
  //: joint g7 (w3) @(289, 322) /w:[ 70 69 72 74 ]
  //: joint g15 (w3) @(289, 163) /w:[ 22 21 24 26 ]
  //: joint g17 (w3) @(289, 113) /w:[ 5 6 12 14 ]
  //: joint g14 (w3) @(289, 183) /w:[ 28 27 30 32 ]
  //: joint g5 (w3) @(289, 363) /w:[ 82 81 84 86 ]
  assign Sa = {w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w3, w2, w3, w3}; //: CONCAT g0  @(352,228) /sn:0 /w:[ 1 89 91 83 85 77 79 71 73 65 67 59 61 53 55 47 49 41 43 35 37 29 31 23 25 17 19 13 0 11 1 3 9 ] /dr:1 /tp:0 /drp:1
  //: joint g18 (w3) @(322, 73) /w:[ 8 -1 7 10 ]
  //: joint g12 (w3) @(289, 224) /w:[ 40 39 42 44 ]

endmodule
//: /netlistEnd

//: /netlistBegin LatchD
module LatchD(Q, D, C, nQ);
//: interface  /sz:(75, 48) /bd:[ Li0>D(14/48) Li1>C(29/48) Ro0<Q(12/48) Ro1<nQ(31/48) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output nQ;    //: /sn:0 {0}(344,179)(388,179){1}
//: {2}(392,179)(416,179)(416,162)(429,162){3}
//: {4}(390,177)(390,132)(300,132)(300,119)(318,119){5}
output Q;    //: /sn:0 {0}(339,117)(379,117){1}
//: {2}(383,117)(425,117)(425,103)(438,103){3}
//: {4}(381,119)(381,161)(313,161)(313,176)(323,176){5}
input C;    //: /sn:0 {0}(25,183)(106,183)(106,160)(138,160){1}
//: {2}(142,160)(181,160){3}
//: {4}(140,158)(140,107)(180,107){5}
input D;    //: /sn:0 {0}(86,90)(118,90){1}
//: {2}(122,90)(167,90)(167,102)(180,102){3}
//: {4}(120,92)(120,155)(181,155){5}
wire w2;    //: /sn:0 {0}(201,105)(303,105)(303,114)(318,114){1}
wire w5;    //: /sn:0 {0}(202,158)(216,158)(216,194)(223,194)(223,181)(323,181){1}
//: enddecls

  //: joint g8 (D) @(120, 90) /w:[ 2 -1 1 4 ]
  //: OUT g4 (Q) @(435,103) /sn:0 /w:[ 3 ]
  _GGNOR2 #(4) g3 (.I0(Q), .I1(w5), .Z(nQ));   //: @(334,179) /sn:0 /w:[ 5 1 0 ]
  _GGNOR2 #(4) g2 (.I0(w2), .I1(nQ), .Z(Q));   //: @(329,117) /sn:0 /w:[ 1 5 0 ]
  _GGAND2 #(6) g1 (.I0(D), .I1(C), .Z(w5));   //: @(192,158) /sn:0 /w:[ 5 3 0 ]
  //: joint g11 (nQ) @(390, 179) /w:[ 2 4 1 -1 ]
  //: joint g10 (Q) @(381, 117) /w:[ 2 -1 1 4 ]
  //: IN g6 (D) @(84,90) /sn:0 /w:[ 0 ]
  //: joint g9 (C) @(140, 160) /w:[ 2 4 1 -1 ]
  //: IN g7 (C) @(23,183) /sn:0 /w:[ 0 ]
  //: OUT g5 (nQ) @(426,162) /sn:0 /w:[ 3 ]
  _GGAND2 #(6) g0 (.I0(!D), .I1(C), .Z(w2));   //: @(191,105) /sn:0 /w:[ 3 5 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin Mux1
module Mux1(Sal, E1, E0, C);
//: interface  /sz:(40, 40) /bd:[ Ti0>C(20/40) Li0>E1(28/40) Li1>E0(10/40) Ro0<Sal(17/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input E1;    //: /sn:0 {0}(293,241)(401,241){1}
input E0;    //: /sn:0 {0}(293,202)(398,202){1}
output Sal;    //: /sn:0 {0}(493,222)(537,222){1}
input C;    //: /sn:0 {0}(359,143)(359,205){1}
//: {2}(361,207)(398,207){3}
//: {4}(359,209)(359,246)(401,246){5}
wire w2;    //: /sn:0 {0}(419,205)(459,205)(459,219)(472,219){1}
wire w5;    //: /sn:0 {0}(422,244)(458,244)(458,224)(472,224){1}
//: enddecls

  _GGAND2 #(6) g4 (.I0(E0), .I1(!C), .Z(w2));   //: @(409,205) /sn:0 /w:[ 1 3 0 ]
  //: OUT g3 (Sal) @(534,222) /sn:0 /w:[ 1 ]
  //: IN g2 (E1) @(291,241) /sn:0 /w:[ 0 ]
  //: IN g1 (E0) @(291,202) /sn:0 /w:[ 0 ]
  _GGOR2 #(6) g6 (.I0(w2), .I1(w5), .Z(Sal));   //: @(483,222) /sn:0 /w:[ 1 1 0 ]
  //: joint g7 (C) @(359, 207) /w:[ 2 1 -1 4 ]
  _GGAND2 #(6) g5 (.I0(E1), .I1(C), .Z(w5));   //: @(412,244) /sn:0 /w:[ 1 5 0 ]
  //: IN g0 (C) @(359,141) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin Mux3x32
module Mux3x32(E0, E2, Sa, E5, E6, E7, E1, E3, C, E4);
//: interface  /sz:(40, 234) /bd:[ Ti0>C[2:0](9/40) Li0>E7[31:0](209/234) Li1>E6[31:0](181/234) Li2>E5[31:0](154/234) Li3>E4[31:0](129/234) Li4>E3[31:0](91/234) Li5>E2[31:0](65/234) Li6>E1[31:0](43/234) Li7>E0[31:0](23/234) Ro0<Sa[31:0](93/234) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [31:0] E7;    //: /sn:0 {0}(#:-80,3036)(-33,3036)(-33,3026)(#:-18,3026){1}
input [31:0] E1;    //: /sn:0 {0}(#:-118,2560)(-33,2560)(-33,2543)(#:-18,2543){1}
output [31:0] Sa;    //: /sn:0 {0}(#:1181,329)(1280,329){1}
input [31:0] E3;    //: /sn:0 {0}(#:-103,2725)(-33,2725)(-33,2704)(#:-18,2704){1}
input [2:0] C;    //: /sn:0 {0}(#:555,-13)(555,-22)(935,-22){1}
//: {2}(937,-24)(#:937,-134){3}
//: {4}(937,-20)(937,129){5}
//: {6}(935,131)(551,131)(#:551,137){7}
//: {8}(937,133)(937,294){9}
//: {10}(935,296)(665,296)(665,274)(551,274)(#:551,284){11}
//: {12}(937,298)(937,406){13}
//: {14}(935,408)(592,408)(592,424)(550,424)(#:550,433){15}
//: {16}(937,410)(937,631){17}
//: {18}(935,633)(605,633)(#:605,641){19}
//: {20}(937,635)(937,786){21}
//: {22}(935,788)(601,788)(#:601,791){23}
//: {24}(937,790)(937,926){25}
//: {26}(935,928)(601,928)(#:601,938){27}
//: {28}(937,930)(937,1071){29}
//: {30}(935,1073)(600,1073)(#:600,1087){31}
//: {32}(937,1075)(937,1259){33}
//: {34}(935,1261)(546,1261)(#:546,1275){35}
//: {36}(937,1263)(937,1410){37}
//: {38}(935,1412)(542,1412)(#:542,1425){39}
//: {40}(937,1414)(937,1569){41}
//: {42}(935,1571)(596,1571)(596,1565)(542,1565)(#:542,1572){43}
//: {44}(937,1573)(937,1700){45}
//: {46}(935,1702)(541,1702)(#:541,1721){47}
//: {48}(937,1704)(937,1956){49}
//: {50}(935,1958)(665,1958)(665,1944)(540,1944)(#:540,1955){51}
//: {52}(937,1960)(937,2101){53}
//: {54}(935,2103)(536,2103)(#:536,2105){55}
//: {56}(937,2105)(937,2247){57}
//: {58}(935,2249)(536,2249)(#:536,2252){59}
//: {60}(937,2251)(937,2377){61}
//: {62}(935,2379)(535,2379)(#:535,2401){63}
//: {64}(937,2381)(937,2633){65}
//: {66}(935,2635)(546,2635)(#:546,2643){67}
//: {68}(937,2637)(937,2786){69}
//: {70}(935,2788)(542,2788)(#:542,2793){71}
//: {72}(937,2790)(937,2946){73}
//: {74}(935,2948)(605,2948)(605,2926)(542,2926)(#:542,2940){75}
//: {76}(937,2950)(937,3073){77}
//: {78}(935,3075)(542,3075)(#:542,3092){79}
//: {80}(937,3077)(937,3253){81}
//: {82}(935,3255)(603,3255)(#:603,3264){83}
//: {84}(937,3257)(937,3407){85}
//: {86}(935,3409)(599,3409)(#:599,3414){87}
//: {88}(937,3411)(937,3553){89}
//: {90}(935,3555)(599,3555)(#:599,3561){91}
//: {92}(937,3557)(937,3699){93}
//: {94}(935,3701)(598,3701)(#:598,3710){95}
//: {96}(937,3703)(937,3995){97}
//: {98}(935,3997)(627,3997)(#:627,4009){99}
//: {100}(937,3999)(937,4155){101}
//: {102}(935,4157)(623,4157)(#:623,4159){103}
//: {104}(937,4159)(937,4302){105}
//: {106}(935,4304)(623,4304)(#:623,4306){107}
//: {108}(937,4306)(937,4436){109}
//: {110}(935,4438)(622,4438)(#:622,4455){111}
//: {112}(937,4440)(937,4726){113}
//: {114}(935,4728)(614,4728)(#:614,4739){115}
//: {116}(937,4730)(937,4879){117}
//: {118}(935,4881)(614,4881)(#:614,4886){119}
//: {120}(937,4883)(937,5025){121}
//: {122}(935,5027)(613,5027)(#:613,5035){123}
//: {124}(937,5029)(937,5180)(613,5180)(#:613,5188){125}
input [31:0] E2;    //: /sn:0 {0}(#:-115,2653)(-33,2653)(-33,2624)(#:-18,2624){1}
input [31:0] E4;    //: /sn:0 {0}(#:-95,2801)(-33,2801)(-33,2784)(#:-18,2784){1}
input [31:0] E6;    //: /sn:0 {0}(#:-89,2954)(-33,2954)(-33,2945)(#:-18,2945){1}
input [31:0] E5;    //: /sn:0 {0}(#:-88,2868)(-33,2868)(-33,2865)(#:-18,2865){1}
input [31:0] E0;    //: /sn:0 {0}(#:-18,2463)(-97,2463)(-97,2462)(#:-121,2462){1}
wire w270;    //: /sn:0 {0}(532,1613)(532,1578){1}
wire w32;    //: /sn:0 {0}(480,257)(520,257){1}
wire w780;    //: /sn:0 {0}(542,5278)(567,5278)(567,5277)(582,5277){1}
wire w341;    //: /sn:0 {0}(504,2481)(464,2481){1}
wire w73;    //: /sn:0 {0}(552,325)(552,305)(551,305)(551,290){1}
wire w405;    //: /sn:0 {0}(511,3001)(486,3001)(486,3000)(471,3000){1}
wire w339;    //: /sn:0 {0}(504,2462)(479,2462)(479,2461)(464,2461){1}
wire w320;    //: /sn:0 {0}(465,2225)(505,2225){1}
wire w244;    //: /sn:0 {0}(470,1831)(510,1831){1}
wire [7:0] w784;    //: /sn:0 {0}(#:536,5273)(39,5273)(39,4955)(#:24,4955){1}
wire w704;    //: /sn:0 {0}(543,4936)(568,4936)(568,4935)(583,4935){1}
wire w699;    //: /sn:0 {0}(646,4389)(673,4389)(673,4254)(805,4254){1}
wire w769;    //: /sn:0 {0}(614,4892)(614,4912)(615,4912)(615,4927){1}
wire w16;    //: /sn:0 {0}(524,48)(499,48)(499,47)(484,47){1}
wire w218;    //: /sn:0 {0}(511,1524)(486,1524)(486,1525)(471,1525){1}
wire w56;    //: /sn:0 {0}(479,503)(504,503)(504,502)(519,502){1}
wire w404;    //: /sn:0 {0}(471,2990)(496,2990)(496,2989)(511,2989){1}
wire w387;    //: /sn:0 {0}(563,2038)(668,2038)(668,2195)(683,2195){1}
wire w4;    //: /sn:0 {0}(524,97)(484,97){1}
wire w616;    //: /sn:0 {0}(592,4239)(552,4239){1}
wire w518;    //: /sn:0 {0}(528,3514)(553,3514)(553,3513)(568,3513){1}
wire w526;    //: /sn:0 {0}(572,3353)(547,3353)(547,3354)(532,3354){1}
wire w628;    //: /sn:0 {0}(556,4119)(596,4119){1}
wire w417;    //: /sn:0 {0}(471,2883)(496,2883)(496,2882)(511,2882){1}
wire w0;    //: /sn:0 {0}(545,-7)(545,28){1}
wire w313;    //: /sn:0 {0}(465,2155)(490,2155)(490,2154)(505,2154){1}
wire w233;    //: /sn:0 {0}(536,1281)(536,1316){1}
wire w240;    //: /sn:0 {0}(470,1791)(495,1791)(495,1790)(510,1790){1}
wire w719;    //: /sn:0 {0}(583,4849)(543,4849){1}
wire w120;    //: /sn:0 {0}(570,911)(530,911){1}
wire w513;    //: /sn:0 {0}(568,3463)(543,3463)(543,3464)(528,3464){1}
wire w641;    //: /sn:0 {0}(591,4535)(551,4535){1}
wire w622;    //: /sn:0 {0}(556,4059)(581,4059)(581,4058)(596,4058){1}
wire w168;    //: /sn:0 {0}(613,979)(613,959)(611,959)(611,944){1}
wire w104;    //: /sn:0 {0}(530,988)(555,988)(555,987)(570,987){1}
wire w111;    //: /sn:0 {0}(530,1058)(570,1058){1}
wire w368;    //: /sn:0 {0}(548,2293)(548,2273)(546,2273)(546,2258){1}
wire w431;    //: /sn:0 {0}(556,2649)(556,2669)(558,2669)(558,2684){1}
wire w287;    //: /sn:0 {0}(569,1358)(678,1358)(678,1519)(693,1519){1}
wire w237;    //: /sn:0 {0}(531,1727)(531,1762){1}
wire w344;    //: /sn:0 {0}(504,2511)(464,2511){1}
wire w119;    //: /sn:0 {0}(530,901)(570,901){1}
wire w54;    //: /sn:0 {0}(479,483)(504,483)(504,482)(519,482){1}
wire w67;    //: /sn:0 {0}(480,374)(505,374)(505,373)(520,373){1}
wire w327;    //: /sn:0 {0}(509,2054)(484,2054)(484,2055)(469,2055){1}
wire w614;    //: /sn:0 {0}(592,4220)(567,4220)(567,4219)(552,4219){1}
wire w745;    //: /sn:0 {0}(582,5155)(542,5155){1}
wire w399;    //: /sn:0 {0}(683,2215)(574,2215)(574,2335)(559,2335){1}
wire w607;    //: /sn:0 {0}(592,4386)(552,4386){1}
wire [7:0] w621;    //: /sn:0 {0}(#:24,4473)(301,4473)(301,4244)(#:546,4244){1}
wire w632;    //: /sn:0 {0}(628,4050)(628,4030)(627,4030)(627,4015){1}
wire [7:0] w167;    //: /sn:0 {0}(#:24,3026)(126,3026)(126,1172)(#:523,1172){1}
wire w587;    //: /sn:0 {0}(744,3507)(737,3507)(737,3347)(626,3347){1}
wire w770;    //: /sn:0 {0}(604,4892)(604,4927){1}
wire w445;    //: /sn:0 {0}(510,3209)(470,3209){1}
wire w124;    //: /sn:0 {0}(574,710)(549,710)(549,711)(534,711){1}
wire w606;    //: /sn:0 {0}(592,4375)(567,4375)(567,4376)(552,4376){1}
wire w687;    //: /sn:0 {0}(650,4092)(775,4092)(775,4234)(805,4234){1}
wire [3:0] w20;    //: /sn:0 {0}(#:811,4249)(1129,4249)(1129,354)(#:1175,354){1}
wire [3:0] w23;    //: /sn:0 {0}(#:699,1534)(1068,1534)(1068,314)(#:1175,314){1}
wire w369;    //: /sn:0 {0}(537,2293)(537,2273)(536,2273)(536,2258){1}
wire w108;    //: /sn:0 {0}(570,1027)(545,1027)(545,1028)(530,1028){1}
wire w508;    //: /sn:0 {0}(528,3651)(553,3651)(553,3650)(568,3650){1}
wire w506;    //: /sn:0 {0}(528,3631)(553,3631)(553,3630)(568,3630){1}
wire w225;    //: /sn:0 {0}(475,1355)(515,1355){1}
wire w507;    //: /sn:0 {0}(568,3641)(528,3641){1}
wire w223;    //: /sn:0 {0}(475,1335)(500,1335)(500,1336)(515,1336){1}
wire w300;    //: /sn:0 {0}(546,2111)(546,2131)(548,2131)(548,2146){1}
wire w126;    //: /sn:0 {0}(574,730)(549,730)(549,731)(534,731){1}
wire w437;    //: /sn:0 {0}(531,3130)(531,3115)(532,3115)(532,3098){1}
wire w125;    //: /sn:0 {0}(534,721)(574,721){1}
wire w8;    //: /sn:0 {0}(484,57)(509,57)(509,56)(524,56){1}
wire w202;    //: /sn:0 {0}(532,1431)(532,1466){1}
wire w669;    //: /sn:0 {0}(623,4312)(623,4332)(624,4332)(624,4347){1}
wire w314;    //: /sn:0 {0}(465,2165)(490,2165)(490,2166)(505,2166){1}
wire [7:0] w71;    //: /sn:0 {0}(#:24,2624)(72,2624)(72,369)(#:474,369){1}
wire w238;    //: /sn:0 {0}(470,1771)(494,1771)(494,1770)(510,1770){1}
wire w520;    //: /sn:0 {0}(528,3534)(568,3534){1}
wire w599;    //: /sn:0 {0}(744,3527)(637,3527)(637,3644)(622,3644){1}
wire w487;    //: /sn:0 {0}(569,2726)(664,2726)(664,2894)(679,2894){1}
wire w400;    //: /sn:0 {0}(552,2799)(552,2819)(554,2819)(554,2834){1}
wire w779;    //: /sn:0 {0}(582,5268)(542,5268){1}
wire w633;    //: /sn:0 {0}(617,4050)(617,4015){1}
wire w211;    //: /sn:0 {0}(511,1692)(471,1692){1}
wire w710;    //: /sn:0 {0}(583,4996)(543,4996){1}
wire w738;    //: /sn:0 {0}(542,5085)(567,5085)(567,5084)(582,5084){1}
wire w742;    //: /sn:0 {0}(542,5125)(567,5125)(567,5124)(582,5124){1}
wire w113;    //: /sn:0 {0}(530,841)(555,841)(555,840)(570,840){1}
wire w345;    //: /sn:0 {0}(464,2521)(504,2521){1}
wire w2;    //: /sn:0 {0}(565,-7)(565,13)(567,13)(567,28){1}
wire w515;    //: /sn:0 {0}(568,3483)(543,3483)(543,3484)(528,3484){1}
wire w433;    //: /sn:0 {0}(536,2649)(536,2684){1}
wire [7:0] w367;    //: /sn:0 {0}(#:24,3669)(221,3669)(221,2486)(#:458,2486){1}
wire w316;    //: /sn:0 {0}(465,2185)(505,2185){1}
wire w115;    //: /sn:0 {0}(570,860)(545,860)(545,861)(530,861){1}
wire w570;    //: /sn:0 {0}(589,3567)(589,3602){1}
wire w458;    //: /sn:0 {0}(679,2904)(580,2904)(580,2876)(565,2876){1}
wire w315;    //: /sn:0 {0}(505,2174)(480,2174)(480,2175)(465,2175){1}
wire w224;    //: /sn:0 {0}(515,1344)(490,1344)(490,1345)(475,1345){1}
wire w10;    //: /sn:0 {0}(484,37)(509,37)(509,36)(524,36){1}
wire w601;    //: /sn:0 {0}(624,4200)(624,4185)(623,4185)(623,4165){1}
wire w469;    //: /sn:0 {0}(542,2946)(542,2966)(543,2966)(543,2981){1}
wire w778;    //: /sn:0 {0}(542,5258)(567,5258)(567,5257)(582,5257){1}
wire w510;    //: /sn:0 {0}(528,3671)(568,3671){1}
wire w438;    //: /sn:0 {0}(470,3139)(495,3139)(495,3138)(510,3138){1}
wire w52;    //: /sn:0 {0}(540,439)(540,474){1}
wire w783;    //: /sn:0 {0}(582,5308)(542,5308){1}
wire w509;    //: /sn:0 {0}(568,3660)(543,3660)(543,3661)(528,3661){1}
wire w142;    //: /sn:0 {0}(569,1176)(544,1176)(544,1177)(529,1177){1}
wire w735;    //: /sn:0 {0}(623,5041)(623,5061)(625,5061)(625,5076){1}
wire [7:0] w330;    //: /sn:0 {0}(#:24,3428)(181,3428)(181,2040)(#:463,2040){1}
wire w50;    //: /sn:0 {0}(560,439)(560,459)(562,459)(562,474){1}
wire w416;    //: /sn:0 {0}(511,2873)(471,2873){1}
wire w406;    //: /sn:0 {0}(471,3010)(496,3010)(496,3009)(511,3009){1}
wire w413;    //: /sn:0 {0}(471,2843)(496,2843)(496,2842)(511,2842){1}
wire w527;    //: /sn:0 {0}(532,3364)(557,3364)(557,3363)(572,3363){1}
wire w432;    //: /sn:0 {0}(546,2649)(546,2669)(547,2669)(547,2684){1}
wire w6;    //: /sn:0 {0}(484,77)(506,77)(506,76)(524,76){1}
wire w744;    //: /sn:0 {0}(542,5145)(582,5145){1}
wire w7;    //: /sn:0 {0}(524,67)(484,67){1}
wire w540;    //: /sn:0 {0}(527,3780)(552,3780)(552,3779)(567,3779){1}
wire w329;    //: /sn:0 {0}(509,2075)(469,2075){1}
wire w99;    //: /sn:0 {0}(707,262)(589,262)(589,367)(574,367){1}
wire w61;    //: /sn:0 {0}(519,553)(479,553){1}
wire w609;    //: /sn:0 {0}(592,4405)(567,4405)(567,4406)(552,4406){1}
wire w441;    //: /sn:0 {0}(470,3169)(510,3169){1}
wire w135;    //: /sn:0 {0}(610,1093)(610,1113)(612,1113)(612,1128){1}
wire w625;    //: /sn:0 {0}(596,4089)(556,4089){1}
wire w216;    //: /sn:0 {0}(511,1505)(471,1505){1}
wire w523;    //: /sn:0 {0}(572,3325)(547,3325)(547,3324)(532,3324){1}
wire w640;    //: /sn:0 {0}(551,4525)(576,4525)(576,4524)(591,4524){1}
wire w531;    //: /sn:0 {0}(615,3305)(615,3285)(613,3285)(613,3270){1}
wire w428;    //: /sn:0 {0}(515,2753)(475,2753){1}
wire w425;    //: /sn:0 {0}(475,2723)(515,2723){1}
wire w106;    //: /sn:0 {0}(530,1008)(555,1008)(555,1007)(570,1007){1}
wire w69;    //: /sn:0 {0}(520,394)(480,394){1}
wire w499;    //: /sn:0 {0}(565,3023)(592,3023)(592,2914)(679,2914){1}
wire w429;    //: /sn:0 {0}(475,2763)(515,2763){1}
wire w304;    //: /sn:0 {0}(465,2302)(490,2302)(490,2301)(505,2301){1}
wire w51;    //: /sn:0 {0}(550,439)(550,459)(551,459)(551,474){1}
wire w207;    //: /sn:0 {0}(471,1652)(511,1652){1}
wire w213;    //: /sn:0 {0}(471,1475)(496,1475)(496,1474)(511,1474){1}
wire w239;    //: /sn:0 {0}(470,1781)(495,1781)(495,1782)(510,1782){1}
wire w718;    //: /sn:0 {0}(543,4839)(568,4839)(568,4838)(583,4838){1}
wire w743;    //: /sn:0 {0}(582,5134)(557,5134)(557,5135)(542,5135){1}
wire w709;    //: /sn:0 {0}(543,4986)(568,4986)(568,4985)(583,4985){1}
wire w66;    //: /sn:0 {0}(480,364)(520,364){1}
wire w299;    //: /sn:0 {0}(693,1539)(581,1539)(581,1655)(565,1655){1}
wire w34;    //: /sn:0 {0}(561,143)(561,163)(563,163)(563,178){1}
wire w326;    //: /sn:0 {0}(469,2045)(494,2045)(494,2044)(509,2044){1}
wire w323;    //: /sn:0 {0}(509,2016)(484,2016)(484,2015)(469,2015){1}
wire w87;    //: /sn:0 {0}(573,516)(692,516)(692,272)(707,272){1}
wire w102;    //: /sn:0 {0}(591,797)(591,832){1}
wire w58;    //: /sn:0 {0}(479,523)(504,523)(504,522)(519,522){1}
wire w781;    //: /sn:0 {0}(582,5287)(557,5287)(557,5288)(542,5288){1}
wire [7:0] w321;    //: /sn:0 {0}(#:24,3508)(201,3508)(201,2190)(#:459,2190){1}
wire w307;    //: /sn:0 {0}(505,2332)(465,2332){1}
wire w28;    //: /sn:0 {0}(520,217)(480,217){1}
wire [7:0] w130;    //: /sn:0 {0}(#:24,2784)(93,2784)(93,726)(#:528,726){1}
wire w629;    //: /sn:0 {0}(596,4129)(556,4129){1}
wire w169;    //: /sn:0 {0}(602,979)(602,959)(601,959)(601,944){1}
wire w435;    //: /sn:0 {0}(553,3130)(553,3113)(552,3113)(552,3098){1}
wire w714;    //: /sn:0 {0}(583,4800)(558,4800)(558,4799)(543,4799){1}
wire w132;    //: /sn:0 {0}(606,682)(606,662)(605,662)(605,647){1}
wire w668;    //: /sn:0 {0}(633,4312)(633,4332)(635,4332)(635,4347){1}
wire w343;    //: /sn:0 {0}(504,2500)(479,2500)(479,2501)(464,2501){1}
wire w511;    //: /sn:0 {0}(568,3681)(528,3681){1}
wire w269;    //: /sn:0 {0}(542,1578)(542,1598)(543,1598)(543,1613){1}
wire w25;    //: /sn:0 {0}(480,187)(505,187)(505,186)(520,186){1}
wire w65;    //: /sn:0 {0}(480,354)(505,354)(505,353)(520,353){1}
wire w210;    //: /sn:0 {0}(511,1682)(471,1682){1}
wire [7:0] w121;    //: /sn:0 {0}(#:24,2865)(103,2865)(103,876)(#:524,876){1}
wire w470;    //: /sn:0 {0}(532,2946)(532,2981){1}
wire w736;    //: /sn:0 {0}(613,5041)(613,5061)(614,5061)(614,5076){1}
wire w308;    //: /sn:0 {0}(465,2342)(490,2342)(490,2341)(505,2341){1}
wire w30;    //: /sn:0 {0}(480,237)(505,237)(505,236)(520,236){1}
wire w217;    //: /sn:0 {0}(471,1515)(496,1515)(496,1514)(511,1514){1}
wire w605;    //: /sn:0 {0}(552,4366)(577,4366)(577,4367)(592,4367){1}
wire w812;    //: /sn:0 {0}(636,5271)(781,5271)(781,4976)(796,4976){1}
wire w758;    //: /sn:0 {0}(637,4822)(781,4822)(781,4946)(796,4946){1}
wire w146;    //: /sn:0 {0}(623,1170)(680,1170)(680,901)(695,901){1}
wire w222;    //: /sn:0 {0}(475,1325)(500,1325)(500,1324)(515,1324){1}
wire w500;    //: /sn:0 {0}(611,3455)(611,3435)(609,3435)(609,3420){1}
wire w713;    //: /sn:0 {0}(543,4789)(568,4789)(568,4788)(583,4788){1}
wire w636;    //: /sn:0 {0}(622,4461)(622,4481)(623,4481)(623,4496){1}
wire w57;    //: /sn:0 {0}(519,513)(479,513){1}
wire w49;    //: /sn:0 {0}(707,252)(589,252)(589,220)(574,220){1}
wire w136;    //: /sn:0 {0}(600,1093)(600,1104)(601,1104)(601,1128){1}
wire w139;    //: /sn:0 {0}(529,1147)(554,1147)(554,1148)(569,1148){1}
wire w318;    //: /sn:0 {0}(465,2205)(490,2205)(490,2204)(505,2204){1}
wire w418;    //: /sn:0 {0}(471,2893)(496,2893)(496,2892)(511,2892){1}
wire w610;    //: /sn:0 {0}(552,4416)(592,4416){1}
wire w105;    //: /sn:0 {0}(570,999)(545,999)(545,998)(530,998){1}
wire w604;    //: /sn:0 {0}(552,4356)(577,4356)(577,4355)(592,4355){1}
wire w505;    //: /sn:0 {0}(568,3622)(543,3622)(543,3621)(528,3621){1}
wire w268;    //: /sn:0 {0}(552,1578)(552,1598)(554,1598)(554,1613){1}
wire w72;    //: /sn:0 {0}(561,290)(561,310)(563,310)(563,325){1}
wire [7:0] w33;    //: /sn:0 {0}(#:24,2543)(67,2543)(67,222)(#:474,222){1}
wire w670;    //: /sn:0 {0}(613,4347)(613,4312){1}
wire w440;    //: /sn:0 {0}(470,3159)(495,3159)(495,3158)(510,3158){1}
wire w107;    //: /sn:0 {0}(530,1018)(570,1018){1}
wire w143;    //: /sn:0 {0}(529,1187)(554,1187)(554,1186)(569,1186){1}
wire w436;    //: /sn:0 {0}(542,3130)(542,3098){1}
wire w536;    //: /sn:0 {0}(599,3751)(599,3731)(598,3731)(598,3716){1}
wire w423;    //: /sn:0 {0}(475,2703)(500,2703)(500,2704)(515,2704){1}
wire w145;    //: /sn:0 {0}(529,1207)(569,1207){1}
wire w219;    //: /sn:0 {0}(471,1535)(511,1535){1}
wire w9;    //: /sn:0 {0}(624,4745)(624,4767)(626,4767)(626,4780){1}
wire w337;    //: /sn:0 {0}(525,2442)(525,2407){1}
wire w201;    //: /sn:0 {0}(542,1431)(542,1451)(543,1451)(543,1466){1}
wire w232;    //: /sn:0 {0}(546,1281)(546,1301)(547,1301)(547,1316){1}
wire w305;    //: /sn:0 {0}(505,2313)(480,2313)(480,2312)(465,2312){1}
wire w55;    //: /sn:0 {0}(519,494)(492,494)(492,493)(479,493){1}
wire [7:0] w430;    //: /sn:0 {0}(#:24,3749)(230,3749)(230,2728)(#:469,2728){1}
wire w613;    //: /sn:0 {0}(552,4209)(577,4209)(577,4208)(592,4208){1}
wire w626;    //: /sn:0 {0}(556,4099)(581,4099)(581,4098)(596,4098){1}
wire w122;    //: /sn:0 {0}(534,691)(559,691)(559,690)(574,690){1}
wire w546;    //: /sn:0 {0}(621,3793)(729,3793)(729,3537)(744,3537){1}
wire w214;    //: /sn:0 {0}(511,1486)(486,1486)(486,1485)(471,1485){1}
wire w220;    //: /sn:0 {0}(511,1545)(471,1545){1}
wire [3:0] w14;    //: /sn:0 {0}(#:750,3522)(1120,3522)(1120,344)(#:1175,344){1}
wire w141;    //: /sn:0 {0}(529,1167)(569,1167){1}
wire w528;    //: /sn:0 {0}(572,3374)(532,3374){1}
wire w643;    //: /sn:0 {0}(591,4554)(566,4554)(566,4555)(551,4555){1}
wire [3:0] w38;    //: /sn:0 {0}(#:713,257)(1165,257)(1165,294)(1175,294){1}
wire w514;    //: /sn:0 {0}(528,3474)(553,3474)(553,3475)(568,3475){1}
wire w426;    //: /sn:0 {0}(515,2732)(490,2732)(490,2733)(475,2733){1}
wire w3;    //: /sn:0 {0}(484,107)(524,107){1}
wire w302;    //: /sn:0 {0}(526,2111)(526,2146){1}
wire w408;    //: /sn:0 {0}(471,3030)(496,3030)(496,3029)(511,3029){1}
wire w127;    //: /sn:0 {0}(534,741)(559,741)(559,740)(574,740){1}
wire w128;    //: /sn:0 {0}(574,751)(534,751){1}
wire w424;    //: /sn:0 {0}(515,2712)(490,2712)(490,2713)(475,2713){1}
wire w133;    //: /sn:0 {0}(595,647)(595,682){1}
wire w635;    //: /sn:0 {0}(632,4461)(632,4481)(634,4481)(634,4496){1}
wire w777;    //: /sn:0 {0}(542,5248)(567,5248)(567,5249)(582,5249){1}
wire w558;    //: /sn:0 {0}(744,3517)(637,3517)(637,3497)(622,3497){1}
wire w204;    //: /sn:0 {0}(511,1621)(486,1621)(486,1622)(471,1622){1}
wire w746;    //: /sn:0 {0}(636,5118)(769,5118)(769,4966)(796,4966){1}
wire w623;    //: /sn:0 {0}(596,4070)(571,4070)(571,4069)(556,4069){1}
wire w502;    //: /sn:0 {0}(589,3455)(589,3420){1}
wire w209;    //: /sn:0 {0}(471,1672)(496,1672)(496,1671)(511,1671){1}
wire w708;    //: /sn:0 {0}(583,4975)(558,4975)(558,4976)(543,4976){1}
wire w701;    //: /sn:0 {0}(615,4780)(615,4759)(614,4759)(614,4745){1}
wire w442;    //: /sn:0 {0}(470,3179)(495,3179)(495,3178)(510,3178){1}
wire w501;    //: /sn:0 {0}(600,3455)(600,3435)(599,3435)(599,3420){1}
wire w504;    //: /sn:0 {0}(528,3611)(553,3611)(553,3610)(568,3610){1}
wire w420;    //: /sn:0 {0}(471,2913)(511,2913){1}
wire w215;    //: /sn:0 {0}(471,1495)(496,1495)(496,1494)(511,1494){1}
wire w706;    //: /sn:0 {0}(543,4956)(568,4956)(568,4955)(583,4955){1}
wire w529;    //: /sn:0 {0}(532,3384)(572,3384){1}
wire w311;    //: /sn:0 {0}(465,2372)(505,2372){1}
wire w524;    //: /sn:0 {0}(532,3334)(557,3334)(557,3333)(572,3333){1}
wire w335;    //: /sn:0 {0}(547,2442)(547,2419)(545,2419)(545,2407){1}
wire w36;    //: /sn:0 {0}(541,143)(541,178){1}
wire w532;    //: /sn:0 {0}(604,3305)(604,3285)(603,3285)(603,3270){1}
wire w631;    //: /sn:0 {0}(637,4015)(637,4030)(639,4030)(639,4050){1}
wire w533;    //: /sn:0 {0}(593,3305)(593,3270){1}
wire w242;    //: /sn:0 {0}(470,1811)(495,1811)(495,1810)(510,1810){1}
wire w740;    //: /sn:0 {0}(542,5105)(567,5105)(567,5104)(582,5104){1}
wire w324;    //: /sn:0 {0}(469,2025)(494,2025)(494,2024)(509,2024){1}
wire w444;    //: /sn:0 {0}(470,3199)(510,3199){1}
wire w419;    //: /sn:0 {0}(511,2903)(471,2903){1}
wire [7:0] w467;    //: /sn:0 {0}(#:24,3990)(246,3990)(246,3174)(#:464,3174){1}
wire w158;    //: /sn:0 {0}(695,881)(639,881)(639,874)(624,874){1}
wire w74;    //: /sn:0 {0}(541,325)(541,290){1}
wire w258;    //: /sn:0 {0}(693,1529)(581,1529)(581,1508)(565,1508){1}
wire w35;    //: /sn:0 {0}(551,143)(551,163)(552,163)(552,178){1}
wire w439;    //: /sn:0 {0}(510,3150)(485,3150)(485,3149)(470,3149){1}
wire w711;    //: /sn:0 {0}(583,5006)(543,5006){1}
wire [7:0] w612;    //: /sn:0 {0}(#:24,4553)(317,4553)(317,4391)(#:546,4391){1}
wire w101;    //: /sn:0 {0}(601,797)(601,817)(602,817)(602,832){1}
wire w332;    //: /sn:0 {0}(540,1961)(540,1981)(541,1981)(541,1996){1}
wire w144;    //: /sn:0 {0}(569,1197)(529,1197){1}
wire w716;    //: /sn:0 {0}(583,4819)(543,4819){1}
wire [3:0] w22;    //: /sn:0 {0}(#:689,2210)(1088,2210)(1088,324)(#:1175,324){1}
wire w741;    //: /sn:0 {0}(582,5115)(542,5115){1}
wire w768;    //: /sn:0 {0}(624,4892)(624,4912)(626,4912)(626,4927){1}
wire w117;    //: /sn:0 {0}(530,881)(555,881)(555,880)(570,880){1}
wire w402;    //: /sn:0 {0}(532,2799)(532,2834){1}
wire w720;    //: /sn:0 {0}(543,4859)(583,4859){1}
wire w228;    //: /sn:0 {0}(515,1385)(475,1385){1}
wire w543;    //: /sn:0 {0}(567,3809)(542,3809)(542,3810)(527,3810){1}
wire w12;    //: /sn:0 {0}(695,871)(680,871)(680,724)(628,724){1}
wire w519;    //: /sn:0 {0}(568,3524)(528,3524){1}
wire w401;    //: /sn:0 {0}(542,2799)(542,2819)(543,2819)(543,2834){1}
wire w309;    //: /sn:0 {0}(505,2351)(480,2351)(480,2352)(465,2352){1}
wire w226;    //: /sn:0 {0}(515,1364)(490,1364)(490,1365)(475,1365){1}
wire w542;    //: /sn:0 {0}(527,3800)(552,3800)(552,3799)(567,3799){1}
wire w301;    //: /sn:0 {0}(536,2111)(536,2131)(537,2131)(537,2146){1}
wire w517;    //: /sn:0 {0}(568,3503)(543,3503)(543,3504)(528,3504){1}
wire w608;    //: /sn:0 {0}(552,4396)(577,4396)(577,4395)(592,4395){1}
wire w200;    //: /sn:0 {0}(552,1431)(552,1451)(554,1451)(554,1466){1}
wire w27;    //: /sn:0 {0}(480,207)(503,207)(503,206)(520,206){1}
wire w715;    //: /sn:0 {0}(543,4809)(568,4809)(568,4808)(583,4808){1}
wire w620;    //: /sn:0 {0}(592,4279)(552,4279){1}
wire w468;    //: /sn:0 {0}(552,2946)(552,2966)(554,2966)(554,2981){1}
wire w138;    //: /sn:0 {0}(529,1137)(554,1137)(554,1136)(569,1136){1}
wire w246;    //: /sn:0 {0}(564,1804)(678,1804)(678,1549)(693,1549){1}
wire w544;    //: /sn:0 {0}(527,3820)(567,3820){1}
wire w411;    //: /sn:0 {0}(511,3060)(471,3060){1}
wire w29;    //: /sn:0 {0}(480,227)(505,227)(505,226)(520,226){1}
wire w231;    //: /sn:0 {0}(556,1281)(556,1301)(558,1301)(558,1316){1}
wire w799;    //: /sn:0 {0}(637,4969)(758,4969)(758,4956)(796,4956){1}
wire w707;    //: /sn:0 {0}(583,4966)(543,4966){1}
wire w443;    //: /sn:0 {0}(510,3188)(485,3188)(485,3189)(470,3189){1}
wire [7:0] w312;    //: /sn:0 {0}(#:24,3588)(213,3588)(213,2337)(#:459,2337){1}
wire w322;    //: /sn:0 {0}(469,2005)(494,2005)(494,2004)(509,2004){1}
wire w370;    //: /sn:0 {0}(526,2293)(526,2258){1}
wire [7:0] w421;    //: /sn:0 {0}(#:24,3830)(238,3830)(238,2878)(#:465,2878){1}
wire w317;    //: /sn:0 {0}(505,2194)(480,2194)(480,2195)(465,2195){1}
wire [7:0] w412;    //: /sn:0 {0}(#:24,3910)(243,3910)(243,3025)(#:465,3025){1}
wire [7:0] w530;    //: /sn:0 {0}(#:24,4071)(249,4071)(249,3349)(#:526,3349){1}
wire w637;    //: /sn:0 {0}(612,4461)(612,4496){1}
wire w645;    //: /sn:0 {0}(551,4575)(591,4575){1}
wire [7:0] w721;    //: /sn:0 {0}(#:24,4714)(522,4714)(522,4824)(#:537,4824){1}
wire w60;    //: /sn:0 {0}(479,543)(519,543){1}
wire [7:0] w112;    //: /sn:0 {0}(#:24,2945)(115,2945)(115,1023)(#:524,1023){1}
wire w336;    //: /sn:0 {0}(536,2442)(536,2422)(535,2422)(535,2407){1}
wire w646;    //: /sn:0 {0}(645,4538)(775,4538)(775,4264)(805,4264){1}
wire w516;    //: /sn:0 {0}(528,3494)(568,3494){1}
wire [3:0] w15;    //: /sn:0 {0}(#:1175,364)(1148,364)(1148,4961)(#:802,4961){1}
wire w618;    //: /sn:0 {0}(592,4258)(567,4258)(567,4259)(552,4259){1}
wire w638;    //: /sn:0 {0}(551,4505)(576,4505)(576,4504)(591,4504){1}
wire w535;    //: /sn:0 {0}(610,3751)(610,3731)(608,3731)(608,3716){1}
wire w414;    //: /sn:0 {0}(511,2854)(486,2854)(486,2853)(471,2853){1}
wire w619;    //: /sn:0 {0}(552,4269)(592,4269){1}
wire w615;    //: /sn:0 {0}(552,4229)(577,4229)(577,4228)(592,4228){1}
wire [7:0] w567;    //: /sn:0 {0}(#:24,4312)(274,4312)(274,3795)(#:521,3795){1}
wire w129;    //: /sn:0 {0}(534,761)(574,761){1}
wire w109;    //: /sn:0 {0}(530,1038)(555,1038)(555,1037)(570,1037){1}
wire w306;    //: /sn:0 {0}(465,2322)(490,2322)(490,2321)(505,2321){1}
wire w229;    //: /sn:0 {0}(475,1395)(515,1395){1}
wire w114;    //: /sn:0 {0}(530,851)(555,851)(555,852)(570,852){1}
wire w331;    //: /sn:0 {0}(550,1961)(550,1981)(552,1981)(552,1996){1}
wire w64;    //: /sn:0 {0}(480,344)(505,344)(505,345)(520,345){1}
wire w539;    //: /sn:0 {0}(567,3771)(542,3771)(542,3770)(527,3770){1}
wire w245;    //: /sn:0 {0}(510,1841)(470,1841){1}
wire [7:0] w267;    //: /sn:0 {0}(#:24,3347)(173,3347)(173,1806)(#:464,1806){1}
wire w63;    //: /sn:0 {0}(480,334)(505,334)(505,333)(520,333){1}
wire w627;    //: /sn:0 {0}(596,4108)(571,4108)(571,4109)(556,4109){1}
wire w644;    //: /sn:0 {0}(591,4565)(551,4565){1}
wire [7:0] w767;    //: /sn:0 {0}(#:536,5120)(418,5120)(418,4875)(#:24,4875){1}
wire w537;    //: /sn:0 {0}(588,3751)(588,3716){1}
wire w236;    //: /sn:0 {0}(541,1727)(541,1747)(542,1747)(542,1762){1}
wire w545;    //: /sn:0 {0}(527,3830)(567,3830){1}
wire [3:0] w21;    //: /sn:0 {0}(#:685,2909)(1097,2909)(1097,334)(#:1175,334){1}
wire w705;    //: /sn:0 {0}(583,4947)(558,4947)(558,4946)(543,4946){1}
wire w333;    //: /sn:0 {0}(530,1961)(530,1996){1}
wire w340;    //: /sn:0 {0}(464,2471)(489,2471)(489,2470)(504,2470){1}
wire w199;    //: /sn:0 {0}(695,891)(639,891)(639,1021)(624,1021){1}
wire [7:0] w712;    //: /sn:0 {0}(#:537,4971)(455,4971)(455,4794)(#:24,4794){1}
wire w617;    //: /sn:0 {0}(552,4249)(577,4249)(577,4248)(592,4248){1}
wire w170;    //: /sn:0 {0}(591,979)(591,944){1}
wire w100;    //: /sn:0 {0}(611,797)(611,817)(613,817)(613,832){1}
wire w31;    //: /sn:0 {0}(480,247)(520,247){1}
wire w600;    //: /sn:0 {0}(635,4200)(635,4180)(633,4180)(633,4165){1}
wire [7:0] w230;    //: /sn:0 {0}(#:24,3106)(133,3106)(133,1360)(#:469,1360){1}
wire w538;    //: /sn:0 {0}(527,3760)(552,3760)(552,3759)(567,3759){1}
wire [7:0] w521;    //: /sn:0 {0}(#:24,4151)(260,4151)(260,3499)(#:522,3499){1}
wire w658;    //: /sn:0 {0}(646,4242)(790,4242)(790,4244)(805,4244){1}
wire [3:0] w24;    //: /sn:0 {0}(#:701,886)(1047,886)(1047,304)(1175,304){1}
wire w358;    //: /sn:0 {0}(683,2205)(574,2205)(574,2188)(559,2188){1}
wire w328;    //: /sn:0 {0}(469,2065)(509,2065){1}
wire w776;    //: /sn:0 {0}(582,5237)(557,5237)(557,5238)(542,5238){1}
wire w1;    //: /sn:0 {0}(555,-7)(555,13)(556,13)(556,28){1}
wire w415;    //: /sn:0 {0}(471,2863)(496,2863)(496,2862)(511,2862){1}
wire w310;    //: /sn:0 {0}(505,2362)(465,2362){1}
wire w235;    //: /sn:0 {0}(551,1727)(551,1747)(553,1747)(553,1762){1}
wire w541;    //: /sn:0 {0}(567,3790)(527,3790){1}
wire w241;    //: /sn:0 {0}(510,1801)(470,1801){1}
wire [7:0] w221;    //: /sn:0 {0}(#:24,3186)(145,3186)(145,1510)(#:465,1510){1}
wire w140;    //: /sn:0 {0}(569,1156)(544,1156)(544,1157)(529,1157){1}
wire w409;    //: /sn:0 {0}(471,3040)(486,3040)(486,3039)(511,3039){1}
wire w346;    //: /sn:0 {0}(558,2484)(668,2484)(668,2225)(683,2225){1}
wire w205;    //: /sn:0 {0}(471,1632)(496,1632)(496,1633)(511,1633){1}
wire w782;    //: /sn:0 {0}(542,5298)(582,5298){1}
wire w522;    //: /sn:0 {0}(532,3314)(557,3314)(557,3313)(572,3313){1}
wire w227;    //: /sn:0 {0}(475,1375)(500,1375)(500,1374)(515,1374){1}
wire w116;    //: /sn:0 {0}(530,871)(570,871){1}
wire w786;    //: /sn:0 {0}(613,5194)(613,5214)(614,5214)(614,5229){1}
wire w243;    //: /sn:0 {0}(510,1820)(485,1820)(485,1821)(470,1821){1}
wire [7:0] w212;    //: /sn:0 {0}(#:24,3267)(165,3267)(165,1657)(#:465,1657){1}
wire [7:0] w18;    //: /sn:0 {0}(#:24,2463)(60,2463)(60,72)(#:478,72){1}
wire w118;    //: /sn:0 {0}(570,890)(545,890)(545,891)(530,891){1}
wire w422;    //: /sn:0 {0}(475,2693)(500,2693)(500,2692)(515,2692){1}
wire w68;    //: /sn:0 {0}(480,384)(505,384)(505,383)(520,383){1}
wire w739;    //: /sn:0 {0}(582,5096)(557,5096)(557,5095)(542,5095){1}
wire w338;    //: /sn:0 {0}(464,2451)(489,2451)(489,2450)(504,2450){1}
wire w702;    //: /sn:0 {0}(604,4780)(604,4745){1}
wire w639;    //: /sn:0 {0}(591,4516)(566,4516)(566,4515)(551,4515){1}
wire w407;    //: /sn:0 {0}(511,3020)(471,3020){1}
wire w123;    //: /sn:0 {0}(534,701)(559,701)(559,702)(574,702){1}
wire w525;    //: /sn:0 {0}(532,3344)(572,3344){1}
wire w59;    //: /sn:0 {0}(519,532)(494,532)(494,533)(479,533){1}
wire w427;    //: /sn:0 {0}(475,2743)(500,2743)(500,2742)(515,2742){1}
wire w568;    //: /sn:0 {0}(609,3567)(609,3587)(611,3587)(611,3602){1}
wire w602;    //: /sn:0 {0}(613,4165)(613,4200){1}
wire [7:0] w62;    //: /sn:0 {0}(#:24,2704)(76,2704)(76,518)(#:473,518){1}
wire w319;    //: /sn:0 {0}(505,2215)(465,2215){1}
wire w787;    //: /sn:0 {0}(603,5194)(603,5229){1}
wire w624;    //: /sn:0 {0}(556,4079)(581,4079)(581,4078)(596,4078){1}
wire w137;    //: /sn:0 {0}(590,1093)(590,1128){1}
wire w11;    //: /sn:0 {0}(578,70)(692,70)(692,242)(707,242){1}
wire w110;    //: /sn:0 {0}(570,1048)(530,1048){1}
wire w70;    //: /sn:0 {0}(480,404)(520,404){1}
wire w717;    //: /sn:0 {0}(583,4828)(558,4828)(558,4829)(543,4829){1}
wire w611;    //: /sn:0 {0}(592,4426)(552,4426){1}
wire w785;    //: /sn:0 {0}(623,5194)(623,5214)(625,5214)(625,5229){1}
wire w206;    //: /sn:0 {0}(511,1641)(486,1641)(486,1642)(471,1642){1}
wire w446;    //: /sn:0 {0}(564,3172)(664,3172)(664,2924)(679,2924){1}
wire w5;    //: /sn:0 {0}(484,87)(509,87)(509,86)(524,86){1}
wire [7:0] w667;    //: /sn:0 {0}(#:24,4634)(326,4634)(326,4540)(#:545,4540){1}
wire w208;    //: /sn:0 {0}(511,1661)(486,1661)(486,1662)(471,1662){1}
wire w642;    //: /sn:0 {0}(551,4545)(576,4545)(576,4544)(591,4544){1}
wire w131;    //: /sn:0 {0}(617,682)(617,662)(615,662)(615,647){1}
wire w410;    //: /sn:0 {0}(471,3050)(511,3050){1}
wire w325;    //: /sn:0 {0}(509,2035)(469,2035){1}
wire [7:0] w512;    //: /sn:0 {0}(#:24,4232)(264,4232)(264,3646)(#:522,3646){1}
wire w342;    //: /sn:0 {0}(464,2491)(489,2491)(489,2490)(504,2490){1}
wire w26;    //: /sn:0 {0}(480,197)(505,197)(505,198)(520,198){1}
wire [7:0] w630;    //: /sn:0 {0}(#:550,4094)(287,4094)(287,4392)(#:24,4392){1}
wire w737;    //: /sn:0 {0}(603,5041)(603,5076){1}
wire w569;    //: /sn:0 {0}(599,3567)(599,3587)(600,3587)(600,3602){1}
//: enddecls

  assign {w36, w35, w34} = C; //: CONCAT g4  @(551,138) /sn:0 /R:1 /w:[ 0 0 0 7 ] /dr:0 /tp:0 /drp:0
  assign {w70, w69, w68, w67, w66, w65, w64, w63} = w71; //: CONCAT g8  @(475,369) /sn:0 /R:2 /w:[ 0 1 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign w21 = {w446, w499, w458, w487}; //: CONCAT g140  @(684,2909) /sn:0 /w:[ 0 1 1 0 1 ] /dr:1 /tp:0 /drp:1
  assign {w111, w110, w109, w108, w107, w106, w105, w104} = w112; //: CONCAT g13  @(525,1023) /sn:0 /R:2 /w:[ 0 1 0 1 0 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w311, w310, w309, w308, w307, w306, w305, w304} = w312; //: CONCAT g37  @(460,2337) /sn:0 /R:2 /w:[ 0 1 1 0 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  Mux3 g55 (.C0(w400), .C1(w401), .C2(w402), .E0(w413), .E1(w414), .E2(w415), .E3(w416), .E4(w417), .E5(w418), .E6(w419), .E7(w420), .Sal(w458));   //: @(512, 2835) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>0 Li2>1 Li3>0 Li4>1 Li5>1 Li6>0 Li7>1 Ro0<1 ]
  assign {w502, w501, w500} = C; //: CONCAT g58  @(599,3415) /sn:0 /R:1 /w:[ 1 1 1 87 ] /dr:0 /tp:0 /drp:0
  assign w20 = {w646, w699, w658, w687}; //: CONCAT g139  @(810,4249) /sn:0 /w:[ 0 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: joint g112 (C) @(937, 2788) /w:[ -1 69 70 72 ]
  assign {w633, w632, w631} = C; //: CONCAT g76  @(627,4010) /sn:0 /R:1 /w:[ 1 1 0 99 ] /dr:0 /tp:0 /drp:0
  //: joint g111 (C) @(937, 2948) /w:[ -1 73 74 76 ]
  assign {w0, w1, w2} = C; //: CONCAT g1  @(555,-12) /sn:0 /R:1 /w:[ 0 0 0 0 ] /dr:0 /tp:0 /drp:0
  assign {w533, w532, w531} = C; //: CONCAT g64  @(603,3265) /sn:0 /R:1 /w:[ 1 1 1 83 ] /dr:0 /tp:0 /drp:0
  Mux3 g11 (.C0(w50), .C1(w51), .C2(w52), .E0(w54), .E1(w55), .E2(w56), .E3(w57), .E4(w58), .E5(w59), .E6(w60), .E7(w61), .Sal(w87));   //: @(520, 475) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>0 Li2>1 Li3>0 Li4>1 Li5>0 Li6>1 Li7>0 Ro0<0 ]
  //: IN g130 (E0) @(-123,2462) /sn:0 /w:[ 1 ]
  //: joint g121 (C) @(937, 1261) /w:[ -1 33 34 36 ]
  assign {w233, w232, w231} = C; //: CONCAT g28  @(546,1276) /sn:0 /R:1 /w:[ 0 0 0 35 ] /dr:0 /tp:0 /drp:0
  assign {w420, w419, w418, w417, w416, w415, w414, w413} = w421; //: CONCAT g50  @(466,2878) /sn:0 /R:2 /w:[ 0 1 0 0 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  //: IN g132 (E2) @(-117,2653) /sn:0 /w:[ 0 ]
  Mux3 g19 (.C0(w100), .C1(w101), .C2(w102), .E0(w113), .E1(w114), .E2(w115), .E3(w116), .E4(w117), .E5(w118), .E6(w119), .E7(w120), .Sal(w158));   //: @(571, 833) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>1 Li2>0 Li3>1 Li4>1 Li5>0 Li6>1 Li7>0 Ro0<1 ]
  //: joint g113 (C) @(937, 2635) /w:[ -1 65 66 68 ]
  //: OUT g146 (Sa) @(1277,329) /sn:0 /w:[ 1 ]
  Mux3 g6 (.C0(w34), .C1(w35), .C2(w36), .E0(w25), .E1(w26), .E2(w27), .E3(w28), .E4(w29), .E5(w30), .E6(w31), .E7(w32), .Sal(w49));   //: @(521, 179) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>1 Li2>1 Li3>0 Li4>1 Li5>1 Li6>1 Li7>1 Ro0<1 ]
  assign {w320, w319, w318, w317, w316, w315, w314, w313} = w321; //: CONCAT g38  @(460,2190) /sn:0 /R:2 /w:[ 0 1 0 1 0 1 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: joint g115 (C) @(937, 2249) /w:[ -1 57 58 60 ]
  assign {w61, w60, w59, w58, w57, w56, w55, w54} = w62; //: CONCAT g7  @(474,518) /sn:0 /R:2 /w:[ 1 0 1 0 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w445, w444, w443, w442, w441, w440, w439, w438} = w467; //: CONCAT g53  @(465,3174) /sn:0 /R:2 /w:[ 1 0 1 0 0 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w629, w628, w627, w626, w625, w624, w623, w622} = w630; //: CONCAT g75  @(551,4094) /sn:0 /R:2 /w:[ 1 0 1 0 1 0 1 0 0 ] /dr:0 /tp:0 /drp:0
  //: IN g135 (E5) @(-90,2868) /sn:0 /w:[ 0 ]
  assign {w170, w169, w168} = C; //: CONCAT g20  @(601,939) /sn:0 /R:1 /w:[ 1 1 1 27 ] /dr:0 /tp:0 /drp:0
  Mux3 g31 (.C0(w200), .C1(w201), .C2(w202), .E0(w213), .E1(w214), .E2(w215), .E3(w216), .E4(w217), .E5(w218), .E6(w219), .E7(w220), .Sal(w258));   //: @(512, 1467) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>0 Li2>1 Li3>0 Li4>1 Li5>0 Li6>1 Li7>0 Ro0<1 ]
  //: joint g124 (C) @(937, 788) /w:[ -1 21 22 24 ]
  assign {w329, w328, w327, w326, w325, w324, w323, w322} = w330; //: CONCAT g39  @(464,2040) /sn:0 /R:2 /w:[ 1 0 1 0 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w570, w569, w568} = C; //: CONCAT g68  @(599,3562) /sn:0 /R:1 /w:[ 0 0 0 91 ] /dr:0 /tp:0 /drp:0
  Mux3 g48 (.C0(w368), .C1(w369), .C2(w370), .E0(w304), .E1(w305), .E2(w306), .E3(w307), .E4(w308), .E5(w309), .E6(w310), .E7(w311), .Sal(w399));   //: @(506, 2294) /sz:(52, 85) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Li0>1 Li1>0 Li2>1 Li3>0 Li4>1 Li5>0 Li6>0 Li7>1 Ro0<1 ]
  assign {w145, w144, w143, w142, w141, w140, w139, w138} = w167; //: CONCAT g17  @(524,1172) /sn:0 /R:2 /w:[ 0 1 0 1 0 1 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w211, w210, w209, w208, w207, w206, w205, w204} = w212; //: CONCAT g25  @(466,1657) /sn:0 /R:2 /w:[ 1 1 0 1 0 1 0 1 1 ] /dr:0 /tp:0 /drp:0
  assign {w245, w244, w243, w242, w241, w240, w239, w238} = w267; //: CONCAT g29  @(465,1806) /sn:0 /R:2 /w:[ 1 0 1 0 1 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w433, w432, w431} = C; //: CONCAT g52  @(546,2644) /sn:0 /R:1 /w:[ 0 0 0 67 ] /dr:0 /tp:0 /drp:0
  //: joint g106 (C) @(937, 3701) /w:[ -1 93 94 96 ]
  //: joint g107 (C) @(937, 3555) /w:[ -1 89 90 92 ]
  Mux3 g83 (.C0(w631), .C1(w632), .C2(w633), .E0(w622), .E1(w623), .E2(w624), .E3(w625), .E4(w626), .E5(w627), .E6(w628), .E7(w629), .Sal(w687));   //: @(597, 4051) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Li0>1 Li1>0 Li2>1 Li3>0 Li4>1 Li5>0 Li6>1 Li7>0 Ro0<0 ]
  //: joint g100 (C) @(937, 4728) /w:[ -1 113 114 116 ]
  assign {w120, w119, w118, w117, w116, w115, w114, w113} = w121; //: CONCAT g14  @(525,876) /sn:0 /R:2 /w:[ 1 0 1 0 0 1 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w370, w369, w368} = C; //: CONCAT g44  @(536,2253) /sn:0 /R:1 /w:[ 1 1 1 59 ] /dr:0 /tp:0 /drp:0
  Mux3 g47 (.C0(w331), .C1(w332), .C2(w333), .E0(w322), .E1(w323), .E2(w324), .E3(w325), .E4(w326), .E5(w327), .E6(w328), .E7(w329), .Sal(w387));   //: @(510, 1997) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>0 Li2>1 Li3>0 Li4>1 Li5>0 Li6>1 Li7>0 Ro0<0 ]
  assign {w670, w669, w668} = C; //: CONCAT g80  @(623,4307) /sn:0 /R:1 /w:[ 1 0 0 107 ] /dr:0 /tp:0 /drp:0
  Mux3cableado g94 (.E7(E7), .E6(E6), .E5(E5), .E4(E4), .E3(E3), .E2(E2), .E1(E1), .E0(E0), .S31(w784), .S30(w767), .S29(w712), .S28(w721), .S27(w667), .S26(w612), .S25(w621), .S24(w630), .S23(w567), .S22(w512), .S21(w521), .S20(w530), .S19(w467), .S18(w412), .S17(w421), .S16(w430), .S15(w367), .S14(w312), .S13(w321), .S12(w330), .S11(w267), .S10(w212), .S9(w221), .S8(w230), .S7(w167), .S6(w112), .S5(w121), .S4(w130), .S3(w62), .S2(w71), .S1(w33), .S0(w18));   //: @(-17, 2383) /sz:(40, 2653) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>1 Li5>1 Li6>1 Li7>0 Ro0<1 Ro1<1 Ro2<1 Ro3<0 Ro4<0 Ro5<0 Ro6<0 Ro7<1 Ro8<0 Ro9<0 Ro10<0 Ro11<0 Ro12<0 Ro13<0 Ro14<0 Ro15<0 Ro16<0 Ro17<0 Ro18<0 Ro19<0 Ro20<0 Ro21<0 Ro22<0 Ro23<0 Ro24<0 Ro25<0 Ro26<0 Ro27<0 Ro28<0 Ro29<0 Ro30<0 Ro31<0 ]
  assign {w137, w136, w135} = C; //: CONCAT g21  @(600,1088) /sn:0 /R:1 /w:[ 0 0 0 31 ] /dr:0 /tp:0 /drp:0
  Mux3 g84 (.C0(w668), .C1(w669), .C2(w670), .E0(w604), .E1(w605), .E2(w606), .E3(w607), .E4(w608), .E5(w609), .E6(w610), .E7(w611), .Sal(w699));   //: @(593, 4348) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>0 Li0>1 Li1>1 Li2>0 Li3>0 Li4>1 Li5>0 Li6>1 Li7>0 Ro0<0 ]
  //: joint g105 (C) @(937, 3997) /w:[ -1 97 98 100 ]
  assign w22 = {w346, w399, w358, w387}; //: CONCAT g141  @(688,2210) /sn:0 /w:[ 0 1 0 0 1 ] /dr:1 /tp:0 /drp:1
  Mux3 g23 (.C0(w131), .C1(w132), .C2(w133), .E0(w122), .E1(w123), .E2(w124), .E3(w125), .E4(w126), .E5(w127), .E6(w128), .E7(w129), .Sal(w12));   //: @(575, 683) /sz:(52, 85) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Li0>1 Li1>1 Li2>0 Li3>1 Li4>0 Li5>1 Li6>0 Li7>1 Ro0<1 ]
  assign {w345, w344, w343, w342, w341, w340, w339, w338} = w367; //: CONCAT g41  @(459,2486) /sn:0 /R:2 /w:[ 0 1 1 0 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w333, w332, w331} = C; //: CONCAT g40  @(540,1956) /sn:0 /R:1 /w:[ 0 0 0 51 ] /dr:0 /tp:0 /drp:0
  Mux3 g54 (.C0(w435), .C1(w436), .C2(w437), .E0(w438), .E1(w439), .E2(w440), .E3(w441), .E4(w442), .E5(w443), .E6(w444), .E7(w445), .Sal(w446));   //: @(511, 3131) /sz:(52, 85) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Li0>1 Li1>0 Li2>1 Li3>1 Li4>1 Li5>0 Li6>1 Li7>0 Ro0<0 ]
  assign {w737, w736, w735} = C; //: CONCAT g93  @(613,5036) /sn:0 /R:1 /w:[ 0 0 0 123 ] /dr:0 /tp:0 /drp:0
  //: joint g116 (C) @(937, 1958) /w:[ -1 49 50 52 ]
  //: joint g123 (C) @(937, 928) /w:[ -1 25 26 28 ]
  Mux3 g0 (.C0(w2), .C1(w1), .C2(w0), .E0(w10), .E1(w16), .E2(w8), .E3(w7), .E4(w6), .E5(w5), .E6(w4), .E7(w3), .Sal(w11));   //: @(525, 29) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>0 Li2>1 Li3>0 Li4>1 Li5>1 Li6>0 Li7>1 Ro0<0 ]
  assign {w220, w219, w218, w217, w216, w215, w214, w213} = w221; //: CONCAT g26  @(466,1510) /sn:0 /R:2 /w:[ 1 0 1 0 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w402, w401, w400} = C; //: CONCAT g46  @(542,2794) /sn:0 /R:1 /w:[ 0 0 0 71 ] /dr:0 /tp:0 /drp:0
  Mux3 g90 (.C0(w735), .C1(w736), .C2(w737), .E0(w738), .E1(w739), .E2(w740), .E3(w741), .E4(w742), .E5(w743), .E6(w744), .E7(w745), .Sal(w746));   //: @(583, 5077) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>0 Li2>1 Li3>0 Li4>1 Li5>0 Li6>1 Li7>0 Ro0<0 ]
  assign {w702, w701, w9} = C; //: CONCAT g82  @(614,4740) /sn:0 /R:1 /w:[ 1 1 0 115 ] /dr:0 /tp:0 /drp:0
  //: IN g136 (E6) @(-91,2954) /sn:0 /w:[ 0 ]
  //: joint g128 (C) @(937, 131) /w:[ -1 5 6 8 ]
  assign {w237, w236, w235} = C; //: CONCAT g33  @(541,1722) /sn:0 /R:1 /w:[ 0 0 0 47 ] /dr:0 /tp:0 /drp:0
  Mux3 g91 (.C0(w9), .C1(w701), .C2(w702), .E0(w713), .E1(w714), .E2(w715), .E3(w716), .E4(w717), .E5(w718), .E6(w719), .E7(w720), .Sal(w758));   //: @(584, 4781) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Li0>1 Li1>0 Li2>1 Li3>0 Li4>0 Li5>1 Li6>0 Li7>1 Ro0<0 ]
  assign {w411, w410, w409, w408, w407, w406, w405, w404} = w412; //: CONCAT g49  @(466,3025) /sn:0 /R:2 /w:[ 1 0 0 0 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  //: IN g137 (E7) @(-82,3036) /sn:0 /w:[ 0 ]
  assign {w511, w510, w509, w508, w507, w506, w505, w504} = w512; //: CONCAT g61  @(523,3646) /sn:0 /R:2 /w:[ 1 0 1 0 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w32, w31, w30, w29, w28, w27, w26, w25} = w33; //: CONCAT g3  @(475,222) /sn:0 /R:2 /w:[ 0 0 0 0 1 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w302, w301, w300} = C; //: CONCAT g34  @(536,2106) /sn:0 /R:1 /w:[ 0 0 0 55 ] /dr:0 /tp:0 /drp:0
  assign {w429, w428, w427, w426, w425, w424, w423, w422} = w430; //: CONCAT g51  @(470,2728) /sn:0 /R:2 /w:[ 0 1 0 1 0 1 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w720, w719, w718, w717, w716, w715, w714, w713} = w721; //: CONCAT g86  @(538,4824) /sn:0 /R:2 /w:[ 0 1 0 1 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w745, w744, w743, w742, w741, w740, w739, w738} = w767; //: CONCAT g89  @(537,5120) /sn:0 /R:2 /w:[ 1 0 1 0 1 0 1 0 0 ] /dr:0 /tp:0 /drp:0
  assign {w3, w4, w5, w6, w7, w8, w16, w10} = w18; //: CONCAT g2  @(479,72) /sn:0 /R:2 /w:[ 0 1 0 0 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w545, w544, w543, w542, w541, w540, w539, w538} = w567; //: CONCAT g65  @(522,3795) /sn:0 /R:2 /w:[ 0 0 1 0 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w645, w644, w643, w642, w641, w640, w639, w638} = w667; //: CONCAT g77  @(546,4540) /sn:0 /R:2 /w:[ 0 1 1 0 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  //: joint g110 (C) @(937, 3075) /w:[ -1 77 78 80 ]
  Mux3 g59 (.C0(w431), .C1(w432), .C2(w433), .E0(w422), .E1(w423), .E2(w424), .E3(w425), .E4(w426), .E5(w427), .E6(w428), .E7(w429), .Sal(w487));   //: @(516, 2685) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>1 Li2>0 Li3>1 Li4>0 Li5>1 Li6>0 Li7>1 Ro0<0 ]
  Mux3 g72 (.C0(w568), .C1(w569), .C2(w570), .E0(w504), .E1(w505), .E2(w506), .E3(w507), .E4(w508), .E5(w509), .E6(w510), .E7(w511), .Sal(w599));   //: @(569, 3603) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>0 Li2>1 Li3>0 Li4>1 Li5>0 Li6>1 Li7>0 Ro0<1 ]
  //: joint g98 (C) @(937, 5027) /w:[ -1 121 122 124 ]
  //: joint g99 (C) @(937, 4881) /w:[ -1 117 118 120 ]
  assign {w133, w132, w131} = C; //: CONCAT g16  @(605,642) /sn:0 /R:1 /w:[ 0 1 1 19 ] /dr:0 /tp:0 /drp:0
  Mux3 g96 (.C0(w768), .C1(w769), .C2(w770), .E0(w704), .E1(w705), .E2(w706), .E3(w707), .E4(w708), .E5(w709), .E6(w710), .E7(w711), .Sal(w799));   //: @(584, 4928) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>0 Li2>1 Li3>0 Li4>0 Li5>1 Li6>0 Li7>0 Ro0<0 ]
  //: joint g103 (C) @(937, 4304) /w:[ -1 105 106 108 ]
  //: joint g122 (C) @(937, 1073) /w:[ -1 29 30 32 ]
  assign {w102, w101, w100} = C; //: CONCAT g10  @(601,792) /sn:0 /R:1 /w:[ 0 0 0 23 ] /dr:0 /tp:0 /drp:0
  Mux3 g78 (.C0(w635), .C1(w636), .C2(w637), .E0(w638), .E1(w639), .E2(w640), .E3(w641), .E4(w642), .E5(w643), .E6(w644), .E7(w645), .Sal(w646));   //: @(592, 4497) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>0 Li2>1 Li3>0 Li4>1 Li5>0 Li6>0 Li7>1 Ro0<0 ]
  assign {w783, w782, w781, w780, w779, w778, w777, w776} = w784; //: CONCAT g87  @(537,5273) /sn:0 /R:2 /w:[ 1 0 1 0 1 0 0 1 0 ] /dr:0 /tp:0 /drp:0
  //: joint g129 (C) @(937, -22) /w:[ -1 2 1 4 ]
  assign {w229, w228, w227, w226, w225, w224, w223, w222} = w230; //: CONCAT g27  @(470,1360) /sn:0 /R:2 /w:[ 0 1 0 1 0 1 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w270, w269, w268} = C; //: CONCAT g32  @(542,1573) /sn:0 /R:1 /w:[ 1 0 0 43 ] /dr:0 /tp:0 /drp:0
  //: joint g102 (C) @(937, 4438) /w:[ -1 109 110 112 ]
  assign w24 = {w146, w199, w158, w12}; //: CONCAT g143  @(700,886) /sn:0 /w:[ 0 1 0 0 0 ] /dr:1 /tp:0 /drp:1
  assign {w537, w536, w535} = C; //: CONCAT g69  @(598,3711) /sn:0 /R:1 /w:[ 1 1 1 95 ] /dr:0 /tp:0 /drp:0
  assign {w74, w73, w72} = C; //: CONCAT g9  @(551,285) /sn:0 /R:1 /w:[ 1 1 0 11 ] /dr:0 /tp:0 /drp:0
  assign {w437, w436, w435} = C; //: CONCAT g57  @(542,3093) /sn:0 /R:1 /w:[ 1 1 1 79 ] /dr:0 /tp:0 /drp:0
  //: joint g119 (C) @(937, 1571) /w:[ -1 41 42 44 ]
  assign w23 = {w246, w299, w258, w287}; //: CONCAT g142  @(698,1534) /sn:0 /w:[ 0 1 0 0 1 ] /dr:1 /tp:0 /drp:1
  assign {w129, w128, w127, w126, w125, w124, w123, w122} = w130; //: CONCAT g15  @(529,726) /sn:0 /R:2 /w:[ 0 1 0 1 0 1 0 0 1 ] /dr:0 /tp:0 /drp:0
  Mux3 g71 (.C0(w531), .C1(w532), .C2(w533), .E0(w522), .E1(w523), .E2(w524), .E3(w525), .E4(w526), .E5(w527), .E6(w528), .E7(w529), .Sal(w587));   //: @(573, 3306) /sz:(52, 85) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Li0>1 Li1>0 Li2>1 Li3>1 Li4>0 Li5>1 Li6>0 Li7>1 Ro0<1 ]
  //: IN g131 (E1) @(-120,2560) /sn:0 /w:[ 0 ]
  Mux3 g67 (.C0(w500), .C1(w501), .C2(w502), .E0(w513), .E1(w514), .E2(w515), .E3(w516), .E4(w517), .E5(w518), .E6(w519), .E7(w520), .Sal(w558));   //: @(569, 3456) /sz:(52, 85) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Li0>0 Li1>1 Li2>0 Li3>1 Li4>0 Li5>1 Li6>0 Li7>1 Ro0<1 ]
  //: joint g127 (C) @(937, 296) /w:[ -1 9 10 12 ]
  Mux3 g43 (.C0(w300), .C1(w301), .C2(w302), .E0(w313), .E1(w314), .E2(w315), .E3(w316), .E4(w317), .E5(w318), .E6(w319), .E7(w320), .Sal(w358));   //: @(506, 2147) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>1 Li2>0 Li3>1 Li4>0 Li5>1 Li6>0 Li7>1 Ro0<1 ]
  assign Sa = {w15, w20, w14, w21, w22, w23, w24, w38}; //: CONCAT g145  @(1180,329) /sn:0 /w:[ 0 0 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign {w520, w519, w518, w517, w516, w515, w514, w513} = w521; //: CONCAT g62  @(523,3499) /sn:0 /R:2 /w:[ 0 1 0 1 0 1 0 1 1 ] /dr:0 /tp:0 /drp:0
  assign {w611, w610, w609, w608, w607, w606, w605, w604} = w612; //: CONCAT g73  @(547,4391) /sn:0 /R:2 /w:[ 1 0 1 0 1 1 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w787, w786, w785} = C; //: CONCAT g88  @(613,5189) /sn:0 /R:1 /w:[ 0 0 0 125 ] /dr:0 /tp:0 /drp:0
  //: joint g104 (C) @(937, 4157) /w:[ -1 101 102 104 ]
  assign w14 = {w546, w599, w558, w587}; //: CONCAT g138  @(749,3522) /sn:0 /w:[ 0 1 0 0 0 ] /dr:1 /tp:0 /drp:1
  Mux3 g42 (.C0(w335), .C1(w336), .C2(w337), .E0(w338), .E1(w339), .E2(w340), .E3(w341), .E4(w342), .E5(w343), .E6(w344), .E7(w345), .Sal(w346));   //: @(505, 2443) /sz:(52, 85) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Li0>1 Li1>0 Li2>1 Li3>0 Li4>1 Li5>0 Li6>0 Li7>1 Ro0<0 ]
  assign {w529, w528, w527, w526, w525, w524, w523, w522} = w530; //: CONCAT g63  @(527,3349) /sn:0 /R:2 /w:[ 0 1 0 1 0 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w620, w619, w618, w617, w616, w615, w614, w613} = w621; //: CONCAT g74  @(547,4244) /sn:0 /R:2 /w:[ 1 0 1 0 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  //: joint g109 (C) @(937, 3255) /w:[ -1 81 82 84 ]
  //: IN g133 (E3) @(-105,2725) /sn:0 /w:[ 0 ]
  assign {w52, w51, w50} = C; //: CONCAT g5  @(550,434) /sn:0 /R:1 /w:[ 0 0 0 15 ] /dr:0 /tp:0 /drp:0
  assign {w470, w469, w468} = C; //: CONCAT g56  @(542,2941) /sn:0 /R:1 /w:[ 0 0 0 75 ] /dr:0 /tp:0 /drp:0
  Mux3 g79 (.C0(w600), .C1(w601), .C2(w602), .E0(w613), .E1(w614), .E2(w615), .E3(w616), .E4(w617), .E5(w618), .E6(w619), .E7(w620), .Sal(w658));   //: @(593, 4201) /sz:(52, 85) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Li0>1 Li1>0 Li2>1 Li3>0 Li4>1 Li5>0 Li6>1 Li7>0 Ro0<0 ]
  Mux3 g95 (.C0(w785), .C1(w786), .C2(w787), .E0(w776), .E1(w777), .E2(w778), .E3(w779), .E4(w780), .E5(w781), .E6(w782), .E7(w783), .Sal(w812));   //: @(583, 5230) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>0 Li1>1 Li2>1 Li3>0 Li4>1 Li5>0 Li6>1 Li7>0 Ro0<0 ]
  //: joint g117 (C) @(937, 2103) /w:[ -1 53 54 56 ]
  Mux3 g24 (.C0(w168), .C1(w169), .C2(w170), .E0(w104), .E1(w105), .E2(w106), .E3(w107), .E4(w108), .E5(w109), .E6(w110), .E7(w111), .Sal(w199));   //: @(571, 980) /sz:(52, 85) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Li0>1 Li1>0 Li2>1 Li3>1 Li4>0 Li5>1 Li6>0 Li7>1 Ro0<1 ]
  Mux3 g36 (.C0(w268), .C1(w269), .C2(w270), .E0(w204), .E1(w205), .E2(w206), .E3(w207), .E4(w208), .E5(w209), .E6(w210), .E7(w211), .Sal(w299));   //: @(512, 1614) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>0 Li0>0 Li1>1 Li2>0 Li3>1 Li4>0 Li5>1 Li6>0 Li7>0 Ro0<1 ]
  assign {w711, w710, w709, w708, w707, w706, w705, w704} = w712; //: CONCAT g85  @(538,4971) /sn:0 /R:2 /w:[ 1 1 0 1 1 0 1 0 0 ] /dr:0 /tp:0 /drp:0
  assign {w770, w769, w768} = C; //: CONCAT g92  @(614,4887) /sn:0 /R:1 /w:[ 0 0 0 119 ] /dr:0 /tp:0 /drp:0
  assign w38 = {w87, w99, w49, w11}; //: CONCAT g144  @(712,257) /sn:0 /w:[ 0 1 0 0 1 ] /dr:1 /tp:0 /drp:1
  //: joint g125 (C) @(937, 633) /w:[ -1 17 18 20 ]
  assign w15 = {w812, w746, w799, w758}; //: CONCAT g101  @(801,4961) /sn:0 /w:[ 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign {w637, w636, w635} = C; //: CONCAT g81  @(622,4456) /sn:0 /R:1 /w:[ 0 0 0 111 ] /dr:0 /tp:0 /drp:0
  Mux3 g60 (.C0(w468), .C1(w469), .C2(w470), .E0(w404), .E1(w405), .E2(w406), .E3(w407), .E4(w408), .E5(w409), .E6(w410), .E7(w411), .Sal(w499));   //: @(512, 2982) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>0 Li2>1 Li3>0 Li4>1 Li5>1 Li6>1 Li7>0 Ro0<0 ]
  //: joint g126 (C) @(937, 408) /w:[ -1 13 14 16 ]
  assign {w602, w601, w600} = C; //: CONCAT g70  @(623,4160) /sn:0 /R:1 /w:[ 0 1 1 103 ] /dr:0 /tp:0 /drp:0
  assign {w337, w336, w335} = C; //: CONCAT g45  @(535,2402) /sn:0 /R:1 /w:[ 1 1 1 63 ] /dr:0 /tp:0 /drp:0
  Mux3 g35 (.C0(w231), .C1(w232), .C2(w233), .E0(w222), .E1(w223), .E2(w224), .E3(w225), .E4(w226), .E5(w227), .E6(w228), .E7(w229), .Sal(w287));   //: @(516, 1317) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>1 Li2>0 Li3>1 Li4>0 Li5>1 Li6>0 Li7>1 Ro0<0 ]
  assign {w202, w201, w200} = C; //: CONCAT g22  @(542,1426) /sn:0 /R:1 /w:[ 0 0 0 39 ] /dr:0 /tp:0 /drp:0
  //: joint g120 (C) @(937, 1412) /w:[ -1 37 38 40 ]
  //: joint g114 (C) @(937, 2379) /w:[ -1 61 62 64 ]
  //: IN g97 (C) @(937,-136) /sn:0 /R:3 /w:[ 3 ]
  Mux3 g66 (.C0(w535), .C1(w536), .C2(w537), .E0(w538), .E1(w539), .E2(w540), .E3(w541), .E4(w542), .E5(w543), .E6(w544), .E7(w545), .Sal(w546));   //: @(568, 3752) /sz:(52, 85) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Li0>1 Li1>0 Li2>1 Li3>0 Li4>1 Li5>0 Li6>1 Li7>1 Ro0<0 ]
  Mux3 g18 (.C0(w135), .C1(w136), .C2(w137), .E0(w138), .E1(w139), .E2(w140), .E3(w141), .E4(w142), .E5(w143), .E6(w144), .E7(w145), .Sal(w146));   //: @(570, 1129) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>1 Li2>0 Li3>1 Li4>0 Li5>1 Li6>0 Li7>1 Ro0<0 ]
  Mux3 g12 (.C0(w72), .C1(w73), .C2(w74), .E0(w63), .E1(w64), .E2(w65), .E3(w66), .E4(w67), .E5(w68), .E6(w69), .E7(w70), .Sal(w99));   //: @(521, 326) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Li0>1 Li1>1 Li2>1 Li3>1 Li4>1 Li5>1 Li6>0 Li7>1 Ro0<1 ]
  //: joint g108 (C) @(937, 3409) /w:[ -1 85 86 88 ]
  Mux3 g30 (.C0(w235), .C1(w236), .C2(w237), .E0(w238), .E1(w239), .E2(w240), .E3(w241), .E4(w242), .E5(w243), .E6(w244), .E7(w245), .Sal(w246));   //: @(511, 1763) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Li0>1 Li1>1 Li2>1 Li3>0 Li4>1 Li5>0 Li6>1 Li7>0 Ro0<0 ]
  //: joint g118 (C) @(937, 1702) /w:[ -1 45 46 48 ]
  //: IN g134 (E4) @(-97,2801) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin ControlALU
module ControlALU(E, ALUOp, Sa);
//: interface  /sz:(88, 40) /bd:[ Ti0>ALUOp[1:0](43/88) Li0>E[5:0](18/40) Ro0<Sa[2:0](18/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
supply0 w24;    //: /sn:0 {0}(457,396)(389,396){1}
//: {2}(387,394)(387,376)(424,376){3}
//: {4}(428,376)(457,376){5}
//: {6}(426,378)(426,386)(457,386){7}
//: {8}(385,396)(235,396)(235,192)(329,192){9}
//: {10}(331,190)(331,158){11}
//: {12}(333,156)(343,156)(343,157)(361,157){13}
//: {14}(331,154)(331,131){15}
//: {16}(333,129)(360,129){17}
//: {18}(331,127)(331,109)(360,109){19}
//: {20}(331,194)(331,205){21}
supply1 w25;    //: /sn:0 {0}(302,67)(302,117){1}
//: {2}(304,119)(360,119){3}
//: {4}(302,121)(302,165){5}
//: {6}(304,167)(361,167){7}
//: {8}(302,169)(302,177)(361,177){9}
output [2:0] Sa;    //: /sn:0 {0}(634,193)(#:554,193){1}
input [1:0] ALUOp;    //: /sn:0 {0}(#:506,78)(532,78)(#:532,137){1}
input [5:0] E;    //: /sn:0 {0}(#:303,265)(#:75,265){1}
wire w7;    //: /sn:0 {0}(309,260)(353,260)(353,255)(368,255){1}
wire [2:0] w4;    //: /sn:0 {0}(#:463,386)(497,386)(497,216)(#:512,216){1}
wire w0;    //: /sn:0 {0}(309,240)(346,240)(346,228)(383,228){1}
wire [2:0] w3;    //: /sn:0 {0}(#:458,253)(481,253)(481,195)(#:512,195){1}
wire w20;    //: /sn:0 {0}(384,255)(436,255)(436,253)(452,253){1}
wire [2:0] w1;    //: /sn:0 {0}(#:366,119)(497,119)(497,154)(#:512,154){1}
wire w18;    //: /sn:0 {0}(404,231)(437,231)(437,243)(452,243){1}
wire w8;    //: /sn:0 {0}(309,270)(336,270)(336,246)(355,246)(355,233)(383,233){1}
wire [2:0] w2;    //: /sn:0 {0}(#:367,167)(493,167)(493,171)(#:512,171){1}
wire w10;    //: /sn:0 {0}(309,290)(324,290){1}
wire w5;    //: /sn:0 {0}(309,250)(345,250)(345,271)(399,271)(399,263)(452,263){1}
wire w9;    //: /sn:0 {0}(309,280)(324,280){1}
//: enddecls

  _GGNBUF #(2) g8 (.I(w7), .Z(w20));   //: @(374,255) /sn:0 /w:[ 1 0 ]
  assign {w10, w9, w8, w7, w5, w0} = E; //: CONCAT g4  @(304,265) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 ] /dr:0 /tp:0 /drp:0
  //: IN g3 (E) @(73,265) /sn:0 /w:[ 1 ]
  //: joint g13 (w25) @(302, 167) /w:[ 6 5 -1 8 ]
  //: IN g2 (ALUOp) @(504,78) /sn:0 /w:[ 0 ]
  //: OUT g1 (Sa) @(631,193) /sn:0 /w:[ 0 ]
  assign w4 = {w24, w24, w24}; //: CONCAT g16  @(462,386) /sn:0 /w:[ 0 0 7 5 ] /dr:1 /tp:0 /drp:1
  //: VDD g11 (w25) @(313,67) /sn:0 /w:[ 0 ]
  //: GROUND g10 (w24) @(331,211) /sn:0 /w:[ 21 ]
  //: joint g19 (w24) @(426, 376) /w:[ 4 -1 3 6 ]
  assign w2 = {w25, w25, w24}; //: CONCAT g6  @(366,167) /sn:0 /w:[ 0 9 7 13 ] /dr:1 /tp:0 /drp:1
  assign w3 = {w5, w20, w18}; //: CONCAT g9  @(457,253) /sn:0 /w:[ 0 1 1 1 ] /dr:1 /tp:0 /drp:1
  _GGOR2 #(6) g7 (.I0(w0), .I1(w8), .Z(w18));   //: @(394,231) /sn:0 /w:[ 1 1 0 ]
  //: joint g15 (w24) @(331, 156) /w:[ 12 14 -1 11 ]
  //: joint g17 (w24) @(331, 192) /w:[ -1 10 9 20 ]
  //: joint g14 (w25) @(302, 119) /w:[ 2 1 -1 4 ]
  assign w1 = {w24, w25, w24}; //: CONCAT g5  @(365,119) /sn:0 /w:[ 0 17 3 19 ] /dr:1 /tp:0 /drp:1
  Mux2x3 g0 (.C(ALUOp), .E3(w4), .E2(w3), .E1(w2), .E0(w1), .Sa(Sa));   //: @(513, 138) /sz:(40, 96) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Li2>1 Li3>1 Ro0<1 ]
  //: joint g18 (w24) @(387, 396) /w:[ 1 2 8 -1 ]
  //: joint g12 (w24) @(331, 129) /w:[ 16 18 -1 15 ]

endmodule
//: /netlistEnd

//: /netlistBegin Mux3cableado
module Mux3cableado(S0, E4, S29, S26, S5, E3, E2, E1, S8, S3, S20, S2, S24, S19, S11, S30, E6, S1, E7, S23, S12, S7, S31, S21, S17, S9, S6, E5, S28, S16, S13, S15, S27, S18, S14, E0, S10, S4, S25, S22);
//: interface  /sz:(40, 2653) /bd:[ Li0>E7[31:0](643/2653) Li1>E6[31:0](562/2653) Li2>E5[31:0](482/2653) Li3>E4[31:0](401/2653) Li4>E3[31:0](321/2653) Li5>E2[31:0](241/2653) Li6>E1[31:0](160/2653) Li7>E0[31:0](80/2653) Ro0<S31[7:0](2572/2653) Ro1<S30[7:0](2492/2653) Ro2<S29[7:0](2411/2653) Ro3<S28[7:0](2331/2653) Ro4<S27[7:0](2251/2653) Ro5<S26[7:0](2170/2653) Ro6<S25[7:0](2090/2653) Ro7<S24[7:0](2009/2653) Ro8<S23[7:0](1929/2653) Ro9<S22[7:0](1849/2653) Ro10<S21[7:0](1768/2653) Ro11<S20[7:0](1688/2653) Ro12<S19[7:0](1607/2653) Ro13<S18[7:0](1527/2653) Ro14<S17[7:0](1447/2653) Ro15<S16[7:0](1366/2653) Ro16<S15[7:0](1286/2653) Ro17<S14[7:0](1205/2653) Ro18<S13[7:0](1125/2653) Ro19<S12[7:0](1045/2653) Ro20<S11[7:0](964/2653) Ro21<S10[7:0](884/2653) Ro22<S9[7:0](803/2653) Ro23<S8[7:0](723/2653) Ro24<S7[7:0](643/2653) Ro25<S6[7:0](562/2653) Ro26<S5[7:0](482/2653) Ro27<S4[7:0](401/2653) Ro28<S3[7:0](321/2653) Ro29<S2[7:0](241/2653) Ro30<S1[7:0](160/2653) Ro31<S0[7:0](80/2653) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [31:0] E7;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [7:0] S7;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E1;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [7:0] S24;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S28;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S13;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E3;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [7:0] S29;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S23;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S2;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S1;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S25;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S12;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E2;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [7:0] S26;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S18;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S27;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S0;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E4;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [7:0] S31;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S10;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E6;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [7:0] S11;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S4;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S8;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S17;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S21;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S20;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S19;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E5;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [7:0] S6;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S16;    //: /sn:0 {0}(#:1,1)(1,1){1}
input [31:0] E0;    //: /sn:0 {0}(#:1,1)(#:1,1){1}
output [7:0] S15;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S9;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S5;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S30;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S14;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S22;    //: /sn:0 {0}(#:1,1)(1,1){1}
output [7:0] S3;    //: /sn:0 {0}(#:1,1)(1,1){1}
wire w32;    //: /sn:0 {0}(1,1)(1,1){1}
wire w73;    //: /sn:0 {0}(1,1)(1,1){1}
wire w45;    //: /sn:0 {0}(1,1)(1,1){1}
wire w96;    //: /sn:0 {0}(1,1)(1,1){1}
wire w160;    //: /sn:0 {0}(1,1)(1,1){1}
wire w244;    //: /sn:0 {0}(1,1)(1,1){1}
wire w218;    //: /sn:0 {0}(1,1)(1,1){1}
wire w56;    //: /sn:0 {0}(1,1)(1,1){1}
wire w16;    //: /sn:0 {0}(1,1)(1,1){1}
wire w81;    //: /sn:0 {0}(1,1)(1,1){1}
wire w19;    //: /sn:0 {0}(1,1)(1,1){1}
wire w4;    //: /sn:0 {0}(1,1)(1,1){1}
wire w89;    //: /sn:0 {0}(1,1)(1,1){1}
wire w183;    //: /sn:0 {0}(1,1)(1,1){1}
wire w0;    //: /sn:0 {0}(1,1)(1,1){1}
wire w151;    //: /sn:0 {0}(1,1)(1,1){1}
wire w240;    //: /sn:0 {0}(1,1)(1,1){1}
wire w233;    //: /sn:0 {0}(1,1)(1,1){1}
wire w120;    //: /sn:0 {0}(1,1)(1,1){1}
wire w104;    //: /sn:0 {0}(1,1)(1,1){1}
wire w111;    //: /sn:0 {0}(1,1)(1,1){1}
wire w168;    //: /sn:0 {0}(1,1)(1,1){1}
wire w171;    //: /sn:0 {0}(1,1)(1,1){1}
wire w237;    //: /sn:0 {0}(1,1)(1,1){1}
wire w67;    //: /sn:0 {0}(1,1)(1,1){1}
wire w54;    //: /sn:0 {0}(1,1)(1,1){1}
wire w119;    //: /sn:0 {0}(1,1)(1,1){1}
wire w90;    //: /sn:0 {0}(1,1)(1,1){1}
wire w176;    //: /sn:0 {0}(1,1)(1,1){1}
wire w167;    //: /sn:0 {0}(1,1)(1,1){1}
wire w23;    //: /sn:0 {0}(1,1)(1,1){1}
wire w20;    //: /sn:0 {0}(1,1)(1,1){1}
wire w124;    //: /sn:0 {0}(1,1)(1,1){1}
wire w174;    //: /sn:0 {0}(1,1)(1,1){1}
wire w225;    //: /sn:0 {0}(1,1)(1,1){1}
wire w108;    //: /sn:0 {0}(1,1)(1,1){1}
wire w223;    //: /sn:0 {0}(1,1)(1,1){1}
wire w126;    //: /sn:0 {0}(1,1)(1,1){1}
wire w125;    //: /sn:0 {0}(1,1)(1,1){1}
wire w8;    //: /sn:0 {0}(1,1)(1,1){1}
wire w103;    //: /sn:0 {0}(1,1)(1,1){1}
wire w238;    //: /sn:0 {0}(1,1)(1,1){1}
wire w71;    //: /sn:0 {0}(1,1)(1,1){1}
wire w202;    //: /sn:0 {0}(1,1)(1,1){1}
wire w17;    //: /sn:0 {0}(1,1)(1,1){1}
wire w84;    //: /sn:0 {0}(1,1)(1,1){1}
wire w53;    //: /sn:0 {0}(1,1)(1,1){1}
wire w255;    //: /sn:0 {0}(1,1)(1,1){1}
wire w211;    //: /sn:0 {0}(1,1)(1,1){1}
wire w44;    //: /sn:0 {0}(1,1)(1,1){1}
wire w2;    //: /sn:0 {0}(1,1)(1,1){1}
wire w113;    //: /sn:0 {0}(1,1)(1,1){1}
wire w83;    //: /sn:0 {0}(1,1)(1,1){1}
wire w77;    //: /sn:0 {0}(1,1)(1,1){1}
wire w115;    //: /sn:0 {0}(1,1)(1,1){1}
wire w224;    //: /sn:0 {0}(1,1)(1,1){1}
wire w10;    //: /sn:0 {0}(1,1)(1,1){1}
wire w190;    //: /sn:0 {0}(1,1)(1,1){1}
wire w52;    //: /sn:0 {0}(1,1)(1,1){1}
wire w95;    //: /sn:0 {0}(1,1)(1,1){1}
wire w188;    //: /sn:0 {0}(1,1)(1,1){1}
wire w142;    //: /sn:0 {0}(1,1)(1,1){1}
wire w155;    //: /sn:0 {0}(1,1)(1,1){1}
wire w178;    //: /sn:0 {0}(1,1)(1,1){1}
wire w187;    //: /sn:0 {0}(1,1)(1,1){1}
wire w50;    //: /sn:0 {0}(1,1)(1,1){1}
wire w6;    //: /sn:0 {0}(1,1)(1,1){1}
wire w7;    //: /sn:0 {0}(1,1)(1,1){1}
wire w93;    //: /sn:0 {0}(1,1)(1,1){1}
wire w61;    //: /sn:0 {0}(1,1)(1,1){1}
wire w99;    //: /sn:0 {0}(1,1)(1,1){1}
wire w135;    //: /sn:0 {0}(1,1)(1,1){1}
wire w153;    //: /sn:0 {0}(1,1)(1,1){1}
wire w216;    //: /sn:0 {0}(1,1)(1,1){1}
wire w239;    //: /sn:0 {0}(1,1)(1,1){1}
wire w69;    //: /sn:0 {0}(1,1)(1,1){1}
wire w51;    //: /sn:0 {0}(1,1)(1,1){1}
wire w106;    //: /sn:0 {0}(1,1)(1,1){1}
wire w207;    //: /sn:0 {0}(1,1)(1,1){1}
wire w213;    //: /sn:0 {0}(1,1)(1,1){1}
wire w66;    //: /sn:0 {0}(1,1)(1,1){1}
wire w37;    //: /sn:0 {0}(1,1)(1,1){1}
wire w177;    //: /sn:0 {0}(1,1)(1,1){1}
wire w234;    //: /sn:0 {0}(1,1)(1,1){1}
wire w34;    //: /sn:0 {0}(1,1)(1,1){1}
wire w254;    //: /sn:0 {0}(1,1)(1,1){1}
wire w87;    //: /sn:0 {0}(1,1)(1,1){1}
wire w43;    //: /sn:0 {0}(1,1)(1,1){1}
wire w102;    //: /sn:0 {0}(1,1)(1,1){1}
wire w157;    //: /sn:0 {0}(1,1)(1,1){1}
wire w58;    //: /sn:0 {0}(1,1)(1,1){1}
wire w28;    //: /sn:0 {0}(1,1)(1,1){1}
wire w130;    //: /sn:0 {0}(1,1)(1,1){1}
wire w169;    //: /sn:0 {0}(1,1)(1,1){1}
wire w132;    //: /sn:0 {0}(1,1)(1,1){1}
wire w184;    //: /sn:0 {0}(1,1)(1,1){1}
wire w25;    //: /sn:0 {0}(1,1)(1,1){1}
wire w65;    //: /sn:0 {0}(1,1)(1,1){1}
wire w210;    //: /sn:0 {0}(1,1)(1,1){1}
wire w40;    //: /sn:0 {0}(1,1)(1,1){1}
wire w92;    //: /sn:0 {0}(1,1)(1,1){1}
wire w121;    //: /sn:0 {0}(1,1)(1,1){1}
wire w217;    //: /sn:0 {0}(1,1)(1,1){1}
wire w30;    //: /sn:0 {0}(1,1)(1,1){1}
wire w162;    //: /sn:0 {0}(1,1)(1,1){1}
wire w222;    //: /sn:0 {0}(1,1)(1,1){1}
wire w146;    //: /sn:0 {0}(1,1)(1,1){1}
wire w149;    //: /sn:0 {0}(1,1)(1,1){1}
wire w165;    //: /sn:0 {0}(1,1)(1,1){1}
wire w248;    //: /sn:0 {0}(1,1)(1,1){1}
wire w57;    //: /sn:0 {0}(1,1)(1,1){1}
wire w49;    //: /sn:0 {0}(1,1)(1,1){1}
wire w136;    //: /sn:0 {0}(1,1)(1,1){1}
wire w139;    //: /sn:0 {0}(1,1)(1,1){1}
wire w173;    //: /sn:0 {0}(1,1)(1,1){1}
wire w252;    //: /sn:0 {0}(1,1)(1,1){1}
wire w105;    //: /sn:0 {0}(1,1)(1,1){1}
wire w148;    //: /sn:0 {0}(1,1)(1,1){1}
wire w186;    //: /sn:0 {0}(1,1)(1,1){1}
wire w72;    //: /sn:0 {0}(1,1)(1,1){1}
wire w94;    //: /sn:0 {0}(1,1)(1,1){1}
wire w33;    //: /sn:0 {0}(1,1)(1,1){1}
wire w191;    //: /sn:0 {0}(1,1)(1,1){1}
wire w107;    //: /sn:0 {0}(1,1)(1,1){1}
wire w143;    //: /sn:0 {0}(1,1)(1,1){1}
wire w219;    //: /sn:0 {0}(1,1)(1,1){1}
wire w79;    //: /sn:0 {0}(1,1)(1,1){1}
wire w9;    //: /sn:0 {0}(1,1)(1,1){1}
wire w145;    //: /sn:0 {0}(1,1)(1,1){1}
wire w232;    //: /sn:0 {0}(1,1)(1,1){1}
wire w55;    //: /sn:0 {0}(1,1)(1,1){1}
wire w39;    //: /sn:0 {0}(1,1)(1,1){1}
wire w201;    //: /sn:0 {0}(1,1)(1,1){1}
wire w122;    //: /sn:0 {0}(1,1)(1,1){1}
wire w134;    //: /sn:0 {0}(1,1)(1,1){1}
wire w166;    //: /sn:0 {0}(1,1)(1,1){1}
wire w203;    //: /sn:0 {0}(1,1)(1,1){1}
wire w214;    //: /sn:0 {0}(1,1)(1,1){1}
wire w220;    //: /sn:0 {0}(1,1)(1,1){1}
wire w14;    //: /sn:0 {0}(1,1)(1,1){1}
wire w141;    //: /sn:0 {0}(1,1)(1,1){1}
wire w179;    //: /sn:0 {0}(1,1)(1,1){1}
wire w250;    //: /sn:0 {0}(1,1)(1,1){1}
wire w38;    //: /sn:0 {0}(1,1)(1,1){1}
wire w195;    //: /sn:0 {0}(1,1)(1,1){1}
wire w152;    //: /sn:0 {0}(1,1)(1,1){1}
wire w180;    //: /sn:0 {0}(1,1)(1,1){1}
wire w182;    //: /sn:0 {0}(1,1)(1,1){1}
wire w3;    //: /sn:0 {0}(1,1)(1,1){1}
wire w181;    //: /sn:0 {0}(1,1)(1,1){1}
wire w194;    //: /sn:0 {0}(1,1)(1,1){1}
wire w127;    //: /sn:0 {0}(1,1)(1,1){1}
wire w128;    //: /sn:0 {0}(1,1)(1,1){1}
wire w133;    //: /sn:0 {0}(1,1)(1,1){1}
wire w75;    //: /sn:0 {0}(1,1)(1,1){1}
wire w204;    //: /sn:0 {0}(1,1)(1,1){1}
wire w209;    //: /sn:0 {0}(1,1)(1,1){1}
wire w215;    //: /sn:0 {0}(1,1)(1,1){1}
wire w156;    //: /sn:0 {0}(1,1)(1,1){1}
wire w41;    //: /sn:0 {0}(1,1)(1,1){1}
wire w36;    //: /sn:0 {0}(1,1)(1,1){1}
wire w242;    //: /sn:0 {0}(1,1)(1,1){1}
wire w82;    //: /sn:0 {0}(1,1)(1,1){1}
wire w74;    //: /sn:0 {0}(1,1)(1,1){1}
wire w158;    //: /sn:0 {0}(1,1)(1,1){1}
wire w35;    //: /sn:0 {0}(1,1)(1,1){1}
wire w91;    //: /sn:0 {0}(1,1)(1,1){1}
wire w101;    //: /sn:0 {0}(1,1)(1,1){1}
wire w163;    //: /sn:0 {0}(1,1)(1,1){1}
wire w192;    //: /sn:0 {0}(1,1)(1,1){1}
wire w22;    //: /sn:0 {0}(1,1)(1,1){1}
wire w144;    //: /sn:0 {0}(1,1)(1,1){1}
wire w117;    //: /sn:0 {0}(1,1)(1,1){1}
wire w172;    //: /sn:0 {0}(1,1)(1,1){1}
wire w228;    //: /sn:0 {0}(1,1)(1,1){1}
wire w12;    //: /sn:0 {0}(1,1)(1,1){1}
wire w226;    //: /sn:0 {0}(1,1)(1,1){1}
wire w78;    //: /sn:0 {0}(1,1)(1,1){1}
wire w200;    //: /sn:0 {0}(1,1)(1,1){1}
wire w27;    //: /sn:0 {0}(1,1)(1,1){1}
wire w246;    //: /sn:0 {0}(1,1)(1,1){1}
wire w86;    //: /sn:0 {0}(1,1)(1,1){1}
wire w138;    //: /sn:0 {0}(1,1)(1,1){1}
wire w231;    //: /sn:0 {0}(1,1)(1,1){1}
wire w80;    //: /sn:0 {0}(1,1)(1,1){1}
wire w29;    //: /sn:0 {0}(1,1)(1,1){1}
wire w42;    //: /sn:0 {0}(1,1)(1,1){1}
wire w147;    //: /sn:0 {0}(1,1)(1,1){1}
wire w247;    //: /sn:0 {0}(1,1)(1,1){1}
wire w60;    //: /sn:0 {0}(1,1)(1,1){1}
wire w46;    //: /sn:0 {0}(1,1)(1,1){1}
wire w112;    //: /sn:0 {0}(1,1)(1,1){1}
wire w175;    //: /sn:0 {0}(1,1)(1,1){1}
wire w15;    //: /sn:0 {0}(1,1)(1,1){1}
wire w109;    //: /sn:0 {0}(1,1)(1,1){1}
wire w129;    //: /sn:0 {0}(1,1)(1,1){1}
wire w229;    //: /sn:0 {0}(1,1)(1,1){1}
wire w97;    //: /sn:0 {0}(1,1)(1,1){1}
wire w114;    //: /sn:0 {0}(1,1)(1,1){1}
wire w245;    //: /sn:0 {0}(1,1)(1,1){1}
wire w64;    //: /sn:0 {0}(1,1)(1,1){1}
wire w63;    //: /sn:0 {0}(1,1)(1,1){1}
wire w159;    //: /sn:0 {0}(1,1)(1,1){1}
wire w236;    //: /sn:0 {0}(1,1)(1,1){1}
wire w76;    //: /sn:0 {0}(1,1)(1,1){1}
wire w21;    //: /sn:0 {0}(1,1)(1,1){1}
wire w170;    //: /sn:0 {0}(1,1)(1,1){1}
wire w199;    //: /sn:0 {0}(1,1)(1,1){1}
wire w249;    //: /sn:0 {0}(1,1)(1,1){1}
wire w230;    //: /sn:0 {0}(1,1)(1,1){1}
wire w31;    //: /sn:0 {0}(1,1)(1,1){1}
wire w100;    //: /sn:0 {0}(1,1)(1,1){1}
wire w251;    //: /sn:0 {0}(1,1)(1,1){1}
wire w24;    //: /sn:0 {0}(1,1)(1,1){1}
wire w1;    //: /sn:0 {0}(1,1)(1,1){1}
wire w161;    //: /sn:0 {0}(1,1)(1,1){1}
wire w241;    //: /sn:0 {0}(1,1)(1,1){1}
wire w235;    //: /sn:0 {0}(1,1)(1,1){1}
wire w221;    //: /sn:0 {0}(1,1)(1,1){1}
wire w140;    //: /sn:0 {0}(1,1)(1,1){1}
wire w196;    //: /sn:0 {0}(1,1)(1,1){1}
wire w253;    //: /sn:0 {0}(1,1)(1,1){1}
wire w154;    //: /sn:0 {0}(1,1)(1,1){1}
wire w205;    //: /sn:0 {0}(1,1)(1,1){1}
wire w227;    //: /sn:0 {0}(1,1)(1,1){1}
wire w98;    //: /sn:0 {0}(1,1)(1,1){1}
wire w116;    //: /sn:0 {0}(1,1)(1,1){1}
wire w243;    //: /sn:0 {0}(1,1)(1,1){1}
wire w18;    //: /sn:0 {0}(1,1)(1,1){1}
wire w118;    //: /sn:0 {0}(1,1)(1,1){1}
wire w212;    //: /sn:0 {0}(1,1)(1,1){1}
wire w68;    //: /sn:0 {0}(1,1)(1,1){1}
wire w164;    //: /sn:0 {0}(1,1)(1,1){1}
wire w198;    //: /sn:0 {0}(1,1)(1,1){1}
wire w59;    //: /sn:0 {0}(1,1)(1,1){1}
wire w123;    //: /sn:0 {0}(1,1)(1,1){1}
wire w85;    //: /sn:0 {0}(1,1)(1,1){1}
wire w62;    //: /sn:0 {0}(1,1)(1,1){1}
wire w185;    //: /sn:0 {0}(1,1)(1,1){1}
wire w11;    //: /sn:0 {0}(1,1)(1,1){1}
wire w137;    //: /sn:0 {0}(1,1)(1,1){1}
wire w197;    //: /sn:0 {0}(1,1)(1,1){1}
wire w70;    //: /sn:0 {0}(1,1)(1,1){1}
wire w110;    //: /sn:0 {0}(1,1)(1,1){1}
wire w150;    //: /sn:0 {0}(1,1)(1,1){1}
wire w189;    //: /sn:0 {0}(1,1)(1,1){1}
wire w193;    //: /sn:0 {0}(1,1)(1,1){1}
wire w206;    //: /sn:0 {0}(1,1)(1,1){1}
wire w88;    //: /sn:0 {0}(1,1)(1,1){1}
wire w13;    //: /sn:0 {0}(1,1)(1,1){1}
wire w48;    //: /sn:0 {0}(1,1)(1,1){1}
wire w5;    //: /sn:0 {0}(1,1)(1,1){1}
wire w208;    //: /sn:0 {0}(1,1)(1,1){1}
wire w47;    //: /sn:0 {0}(1,1)(1,1){1}
wire w131;    //: /sn:0 {0}(1,1)(1,1){1}
wire w26;    //: /sn:0 {0}(1,1)(1,1){1}
//: enddecls

  //: OUT g8 (S0) @(1,1) /sn:0 /w:[ 1 ]
  //: IN g4 (E4) @(1,1) /sn:0 /w:[ 0 ]
  assign S13 = {w237, w205, w173, w141, w109, w77, w45, w13}; //: CONCAT g61  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g37 (S29) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g34 (S26) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g13 (S5) @(1,1) /sn:0 /w:[ 1 ]
  //: IN g3 (E3) @(1,1) /sn:0 /w:[ 0 ]
  assign S10 = {w234, w202, w170, w138, w106, w74, w42, w10}; //: CONCAT g58  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S7 = {w231, w199, w167, w135, w103, w71, w39, w7}; //: CONCAT g55  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S3 = {w227, w195, w163, w131, w99, w67, w35, w3}; //: CONCAT g51  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g2 (E2) @(1,1) /sn:0 /w:[ 0 ]
  assign S29 = {w253, w221, w189, w157, w125, w93, w61, w29}; //: CONCAT g77  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S28 = {w252, w220, w188, w156, w124, w92, w60, w28}; //: CONCAT g76  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S17 = {w241, w209, w177, w145, w113, w81, w49, w17}; //: CONCAT g65  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S11 = {w235, w203, w171, w139, w107, w75, w43, w11}; //: CONCAT g59  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g1 (E1) @(1,1) /sn:0 /w:[ 0 ]
  assign S24 = {w248, w216, w184, w152, w120, w88, w56, w24}; //: CONCAT g72  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S16 = {w240, w208, w176, w144, w112, w80, w48, w16}; //: CONCAT g64  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g16 (S8) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g11 (S3) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g28 (S20) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g10 (S2) @(1,1) /sn:0 /w:[ 1 ]
  assign S30 = {w254, w222, w190, w158, w126, w94, w62, w30}; //: CONCAT g78  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S2 = {w226, w194, w162, w130, w98, w66, w34, w2}; //: CONCAT g50  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g32 (S24) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g27 (S19) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g19 (S11) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g38 (S30) @(1,1) /sn:0 /w:[ 1 ]
  //: IN g6 (E6) @(1,1) /sn:0 /w:[ 0 ]
  assign S21 = {w245, w213, w181, w149, w117, w85, w53, w21}; //: CONCAT g69  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g9 (S1) @(1,1) /sn:0 /w:[ 1 ]
  //: IN g7 (E7) @(1,1) /sn:0 /w:[ 0 ]
  assign S27 = {w251, w219, w187, w155, w123, w91, w59, w27}; //: CONCAT g75  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S9 = {w233, w201, w169, w137, w105, w73, w41, w9}; //: CONCAT g57  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S5 = {w229, w197, w165, w133, w101, w69, w37, w5}; //: CONCAT g53  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g31 (S23) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g20 (S12) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g15 (S7) @(1,1) /sn:0 /w:[ 1 ]
  assign S23 = {w247, w215, w183, w151, w119, w87, w55, w23}; //: CONCAT g71  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g39 (S31) @(1,1) /sn:0 /w:[ 1 ]
  assign S20 = {w244, w212, w180, w148, w116, w84, w52, w20}; //: CONCAT g68  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S19 = {w243, w211, w179, w147, w115, w83, w51, w19}; //: CONCAT g67  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S0 = {w224, w192, w160, w128, w96, w64, w32, w0}; //: CONCAT g48  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign {w127, w126, w125, w124, w123, w122, w121, w120, w119, w118, w117, w116, w115, w114, w113, w112, w111, w110, w109, w108, w107, w106, w105, w104, w103, w102, w101, w100, w99, w98, w97, w96} = E3; //: CONCAT g43  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: OUT g29 (S21) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g25 (S17) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g17 (S9) @(1,1) /sn:0 /w:[ 1 ]
  assign S25 = {w249, w217, w185, w153, w121, w89, w57, w25}; //: CONCAT g73  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S14 = {w238, w206, w174, w142, w110, w78, w46, w14}; //: CONCAT g62  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S15 = {w239, w207, w175, w143, w111, w79, w47, w15}; //: CONCAT g63  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S4 = {w228, w196, w164, w132, w100, w68, w36, w4}; //: CONCAT g52  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign {w95, w94, w93, w92, w91, w90, w89, w88, w87, w86, w85, w84, w83, w82, w81, w80, w79, w78, w77, w76, w75, w74, w73, w72, w71, w70, w69, w68, w67, w66, w65, w64} = E2; //: CONCAT g42  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S26 = {w250, w218, w186, w154, w122, w90, w58, w26}; //: CONCAT g74  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g14 (S6) @(1,1) /sn:0 /w:[ 1 ]
  //: IN g5 (E5) @(1,1) /sn:0 /w:[ 0 ]
  assign S8 = {w232, w200, w168, w136, w104, w72, w40, w8}; //: CONCAT g56  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S31 = {w255, w223, w191, w159, w127, w95, w63, w31}; //: CONCAT g79  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign {w255, w254, w253, w252, w251, w250, w249, w248, w247, w246, w245, w244, w243, w242, w241, w240, w239, w238, w237, w236, w235, w234, w233, w232, w231, w230, w229, w228, w227, w226, w225, w224} = E7; //: CONCAT g47  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w159, w158, w157, w156, w155, w154, w153, w152, w151, w150, w149, w148, w147, w146, w145, w144, w143, w142, w141, w140, w139, w138, w137, w136, w135, w134, w133, w132, w131, w130, w129, w128} = E4; //: CONCAT g44  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: OUT g36 (S28) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g24 (S16) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g21 (S13) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g23 (S15) @(1,1) /sn:0 /w:[ 1 ]
  assign {w63, w62, w61, w60, w59, w58, w57, w56, w55, w54, w53, w52, w51, w50, w49, w48, w47, w46, w45, w44, w43, w42, w41, w40, w39, w38, w37, w36, w35, w34, w33, w32} = E1; //: CONCAT g41  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S12 = {w236, w204, w172, w140, w108, w76, w44, w12}; //: CONCAT g60  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign S6 = {w230, w198, w166, w134, w102, w70, w38, w6}; //: CONCAT g54  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign {w31, w30, w29, w28, w27, w26, w25, w24, w23, w22, w21, w20, w19, w18, w17, w16, w15, w14, w13, w12, w11, w10, w9, w8, w7, w6, w5, w4, w3, w2, w1, w0} = E0; //: CONCAT g40  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: OUT g35 (S27) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g26 (S18) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g22 (S14) @(1,1) /sn:0 /w:[ 1 ]
  //: IN g0 (E0) @(1,1) /sn:0 /w:[ 0 ]
  assign S22 = {w246, w214, w182, w150, w118, w86, w54, w22}; //: CONCAT g70  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign {w223, w222, w221, w220, w219, w218, w217, w216, w215, w214, w213, w212, w211, w210, w209, w208, w207, w206, w205, w204, w203, w202, w201, w200, w199, w198, w197, w196, w195, w194, w193, w192} = E6; //: CONCAT g46  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w191, w190, w189, w188, w187, w186, w185, w184, w183, w182, w181, w180, w179, w178, w177, w176, w175, w174, w173, w172, w171, w170, w169, w168, w167, w166, w165, w164, w163, w162, w161, w160} = E5; //: CONCAT g45  @(1,1) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign S18 = {w242, w210, w178, w146, w114, w82, w50, w18}; //: CONCAT g66  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g18 (S10) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g12 (S4) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g33 (S25) @(1,1) /sn:0 /w:[ 1 ]
  //: OUT g30 (S22) @(1,1) /sn:0 /w:[ 1 ]
  assign S1 = {w225, w193, w161, w129, w97, w65, w33, w1}; //: CONCAT g49  @(1,1) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1

endmodule
//: /netlistEnd

//: /netlistBegin FlipFlopJK
module FlipFlopJK(Q, nQ, J, Reloj, R, K);
//: interface  /sz:(77, 58) /bd:[ Ti0>R(36/77) Li0>J(13/58) Li1>K(39/58) Bi0>Reloj(37/77) Ro0<Q(13/58) Ro1<nQ(39/58) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output Q;    //: /sn:0 {0}(504,284)(531,284){1}
//: {2}(535,284)(551,284)(551,268)(581,268){3}
//: {4}(533,282)(533,173)(184,173)(184,210){5}
//: {6}(186,212)(207,212){7}
//: {8}(184,214)(184,259)(207,259){9}
output nQ;    //: /sn:0 {0}(504,311)(538,311)(538,326)(549,326)(549,342)(581,342){1}
input K;    //: /sn:0 {0}(39,256)(95,256){1}
input R;    //: /sn:0 {0}(70,149)(70,202){1}
//: {2}(72,204)(95,204){3}
//: {4}(70,206)(70,251)(95,251){5}
input J;    //: /sn:0 {0}(95,209)(35,209){1}
supply0 w8;    //: /sn:0 {0}(645,307)(645,241){1}
//: {2}(645,237)(645,220)(653,220){3}
//: {4}(657,220)(673,220){5}
//: {6}(675,218)(675,134)(701,134){7}
//: {8}(675,222)(675,251)(690,251){9}
//: {10}(655,222)(655,256)(690,256){11}
//: {12}(643,239)(631,239)(631,129)(701,129){13}
supply1 w12;    //: /sn:0 {0}(513,367)(513,382)(445,382)(445,336){1}
input Reloj;    //: /sn:0 {0}(228,370)(364,370)(364,308)(373,308){1}
wire w6;    //: /sn:0 {0}(711,256)(813,256)(813,241)(828,241){1}
wire w7;    //: /sn:0 {0}(294,232)(358,232)(358,282)(373,282){1}
wire w14;    //: /sn:0 {0}(228,257)(258,257)(258,234)(273,234){1}
wire w4;    //: /sn:0 {0}(690,261)(680,261)(680,291)(903,291)(903,239)(892,239)(892,238)(886,238){1}
//: {2}(884,236)(884,170)(819,170)(819,156)(831,156){3}
//: {4}(882,238)(864,238)(864,239)(849,239){5}
wire w3;    //: /sn:0 {0}(852,154)(883,154)(883,155)(909,155){1}
//: {2}(911,153)(911,100)(697,100)(697,124)(701,124){3}
//: {4}(911,157)(911,222)(824,222)(824,236)(828,236){5}
wire w2;    //: /sn:0 {0}(722,129)(816,129)(816,151)(831,151){1}
wire w10;    //: /sn:0 {0}(228,210)(258,210)(258,229)(273,229){1}
wire w13;    //: /sn:0 {0}(116,254)(207,254){1}
wire w5;    //: /sn:0 {0}(116,207)(207,207){1}
//: enddecls

  _GGNOR2 #(4) g8 (.I0(w3), .I1(w6), .Z(w4));   //: @(839,239) /sn:0 /w:[ 5 1 5 ]
  //: OUT g4 (Q) @(578,268) /sn:0 /w:[ 3 ]
  //: comment g13 @(640,194) /sn:0
  //: /line:"Reloj"
  //: /end
  //: OUT g3 (nQ) @(578,342) /sn:0 /w:[ 1 ]
  _GGOR2 #(6) g34 (.I0(R), .I1(K), .Z(w13));   //: @(106,254) /sn:0 /w:[ 5 1 0 ]
  //: comment g37 @(89,170) /sn:0
  //: /line:"Reset"
  //: /end
  //: IN g2 (J) @(33,209) /sn:0 /w:[ 1 ]
  //: IN g1 (Reloj) @(226,370) /sn:0 /w:[ 0 ]
  //: comment g16 @(906,244) /sn:0
  //: /line:"nQ"
  //: /end
  //: joint g11 (w4) @(884, 238) /w:[ 1 2 4 -1 ]
  //: joint g10 (w3) @(911, 155) /w:[ -1 2 1 4 ]
  //: joint g28 (w8) @(675, 220) /w:[ -1 6 5 8 ]
  //: VDD g19 (w12) @(524,367) /sn:0 /w:[ 0 ]
  //: GROUND g27 (w8) @(645,313) /sn:0 /w:[ 0 ]
  //: IN g32 (R) @(70,147) /sn:0 /R:3 /w:[ 0 ]
  _GGAND3 #(8) g6 (.I0(w8), .I1(w8), .I2(w4), .Z(w6));   //: @(701,256) /sn:0 /w:[ 9 11 0 0 ]
  //: frame g9 @(625,45) /sn:0 /wi:337 /ht:293 /tx:""
  _GGNOR2 #(4) g7 (.I0(w2), .I1(w4), .Z(w3));   //: @(842,154) /sn:0 /w:[ 1 3 0 ]
  //: comment g15 @(661,256) /sn:0
  //: /line:"J"
  //: /end
  _GGAND2 #(6) g20 (.I0(w5), .I1(!Q), .Z(w10));   //: @(218,210) /sn:0 /w:[ 1 7 0 ]
  //: comment g31 @(374,67) /sn:0
  //: /line:"Flanco ascendente"
  //: /line:""
  //: /line:"Para iniciar poner k a 1 y J a 0"
  //: /line:"Se inicia a 0"
  //: /line:""
  //: /line:"Con poner 1 en R basta"
  //: /end
  //: comment g17 @(917,149) /sn:0
  //: /line:"Q"
  //: /end
  //: frame g25 @(156,145) /sn:0 /wi:159 /ht:135 /tx:""
  //: joint g29 (w8) @(655, 220) /w:[ 4 -1 3 10 ]
  //: comment g14 @(678,114) /sn:0
  //: /line:"K"
  //: /end
  _GGAND3 #(8) g5 (.I0(w3), .I1(w8), .I2(w8), .Z(w2));   //: @(712,129) /sn:0 /w:[ 3 13 7 0 ]
  _GGAND2 #(6) g21 (.I0(!w13), .I1(Q), .Z(w14));   //: @(218,257) /sn:0 /w:[ 1 9 0 ]
  //: joint g24 (Q) @(184, 212) /w:[ 6 5 -1 8 ]
  //: frame g36 @(55,168) /sn:0 /wi:93 /ht:101 /tx:""
  //: joint g23 (Q) @(533, 284) /w:[ 2 4 1 -1 ]
  //: IN g0 (K) @(37,256) /sn:0 /w:[ 0 ]
  _GGOR2 #(6) g22 (.I0(w10), .I1(w14), .Z(w7));   //: @(284,232) /sn:0 /w:[ 1 1 0 ]
  //: comment g26 @(201,148) /sn:0
  //: /line:"Transicion JK"
  //: /end
  //: joint g35 (R) @(70, 204) /w:[ 2 1 -1 4 ]
  FlipFlopD g18 (.Reloj(Reloj), .D(w7), .W(w12), .nQ(nQ), .Q(Q));   //: @(374, 257) /sz:(129, 78) /sn:0 /p:[ Li0>1 Li1>1 Bi0>1 Ro0<0 Ro1<0 ]
  //: comment g12 @(720,56) /sn:0
  //: /line:"Como pone en internet(no funciona)"
  //: /end
  //: joint g30 (w8) @(645, 239) /w:[ -1 2 12 1 ]
  _GGAND2 #(6) g33 (.I0(!R), .I1(J), .Z(w5));   //: @(106,207) /sn:0 /w:[ 3 0 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin ALU1bit
module ALU1bit(B, A, C, AcarreoS, AcarreoE, Sa);
//: interface  /sz:(87, 60) /bd:[ Ti0>AcarreoE(31/87) Ti1>C[2:0](66/87) Li0>A(21/60) Li1>B(36/60) Bo0<AcarreoS(32/87) Ro0<Sa(31/60) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(319,334)(276,334)(276,333)(246,333){1}
//: {2}(242,333)(211,333)(211,332)(203,332){3}
//: {4}(201,330)(201,163)(461,163){5}
//: {6}(465,163)(502,163){7}
//: {8}(463,165)(463,182)(503,182){9}
//: {10}(201,334)(201,379)(88,379){11}
//: {12}(244,335)(244,352)(260,352){13}
input A;    //: /sn:0 {0}(420,245)(407,245)(407,160){1}
//: {2}(409,158)(479,158){3}
//: {4}(483,158)(502,158){5}
//: {6}(481,160)(481,177)(503,177){7}
//: {8}(405,158)(186,158)(186,157)(80,157){9}
input AcarreoE;    //: /sn:0 {0}(433,56)(433,214)(454,214)(454,229){1}
output Sa;    //: /sn:0 {0}(716,201)(901,201)(901,199)(916,199){1}
output AcarreoS;    //: /sn:0 {0}(454,291)(454,348)(465,348)(465,363){1}
supply0 w2;    //: /sn:0 {0}(662,207)(593,207){1}
//: {2}(591,205)(591,198)(662,198){3}
//: {4}(589,207)(579,207)(579,217)(662,217){5}
//: {6}(591,209)(591,236){7}
//: {8}(593,238)(662,238){9}
//: {10}(591,240)(591,264){11}
input [2:0] C;    //: /sn:0 {0}(#:694,69)(#:694,35){1}
wire w6;    //: /sn:0 {0}(523,161)(647,161)(647,167)(662,167){1}
wire w7;    //: /sn:0 {0}(524,180)(647,180)(647,179)(662,179){1}
wire w16;    //: /sn:0 {0}(361,341)(406,341)(406,267)(420,267){1}
wire w0;    //: /sn:0 {0}(704,75)(704,144)(705,144)(705,159){1}
wire w3;    //: /sn:0 {0}(340,323)(340,120)(682,120){1}
//: {2}(684,118)(684,75){3}
//: {4}(684,122)(684,146)(683,146)(683,159){5}
wire w1;    //: /sn:0 {0}(694,75)(694,159){1}
wire w8;    //: /sn:0 {0}(662,228)(555,228)(555,230)(545,230){1}
//: {2}(543,228)(543,187)(662,187){3}
//: {4}(543,232)(543,258)(489,258){5}
wire w22;    //: /sn:0 {0}(276,352)(319,352){1}
//: enddecls

  //: IN g4 (B) @(86,379) /sn:0 /w:[ 11 ]
  Mux3 g8 (.C2(w3), .C1(w1), .C0(w0), .E7(w2), .E6(w8), .E5(w2), .E4(w2), .E3(w2), .E2(w8), .E1(w7), .E0(w6), .Sal(Sa));   //: @(663, 160) /sz:(52, 85) /sn:0 /p:[ Ti0>5 Ti1>1 Ti2>1 Li0>9 Li1>0 Li2>5 Li3>0 Li4>3 Li5>3 Li6>1 Li7>1 Ro0<0 ]
  //: IN g3 (A) @(78,157) /sn:0 /w:[ 9 ]
  //: joint g13 (w8) @(543, 230) /w:[ 1 2 -1 4 ]
  //: GROUND g2 (w2) @(591,270) /sn:0 /w:[ 11 ]
  //: IN g1 (C) @(694,33) /sn:0 /R:3 /w:[ 1 ]
  _GGAND2 #(6) g11 (.I0(A), .I1(B), .Z(w6));   //: @(513,161) /sn:0 /w:[ 5 7 0 ]
  //: joint g16 (A) @(407, 158) /w:[ 2 -1 8 1 ]
  Mux1 g10 (.C(w3), .E1(w22), .E0(B), .Sal(w16));   //: @(320, 324) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Li0>1 Li1>0 Ro0<0 ]
  //: joint g19 (B) @(244, 333) /w:[ 1 -1 2 12 ]
  //: OUT g6 (AcarreoS) @(465,360) /sn:0 /R:3 /w:[ 1 ]
  assign {w3, w1, w0} = C; //: CONCAT g7  @(694,70) /sn:0 /R:1 /w:[ 3 0 0 0 ] /dr:0 /tp:0 /drp:0
  Suma g9 (.AcarreoE(AcarreoE), .A(A), .B(w16), .AcarreoS(AcarreoS), .Suma(w8));   //: @(421, 230) /sz:(67, 60) /sn:0 /p:[ Ti0>1 Li0>0 Li1>1 Bo0<0 Ro0<5 ]
  //: joint g15 (B) @(463, 163) /w:[ 6 -1 5 8 ]
  //: joint g20 (w3) @(684, 120) /w:[ -1 2 1 4 ]
  //: joint g17 (B) @(201, 332) /w:[ 3 4 -1 10 ]
  //: IN g5 (AcarreoE) @(433,54) /sn:0 /R:3 /w:[ 0 ]
  //: joint g14 (A) @(481, 158) /w:[ 4 -1 3 6 ]
  //: joint g21 (w2) @(591, 238) /w:[ 8 7 -1 10 ]
  //: OUT g0 (Sa) @(913,199) /sn:0 /w:[ 1 ]
  //: joint g22 (w2) @(591, 207) /w:[ 1 2 4 6 ]
  _GGOR2 #(6) g12 (.I0(A), .I1(B), .Z(w7));   //: @(514,180) /sn:0 /w:[ 7 9 0 ]
  _GGNBUF #(2) g18 (.I(B), .Z(w22));   //: @(266,352) /sn:0 /w:[ 13 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin Suma
module Suma(AcarreoE, B, Suma, AcarreoS, A);
//: interface  /sz:(67, 60) /bd:[ Ti0>AcarreoE(33/67) Li0>A(15/60) Li1>B(37/60) Bo0<AcarreoS(33/67) Ro0<Suma(28/60) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(98,198)(220,198){1}
//: {2}(224,198)(254,198){3}
//: {4}(258,198)(374,198){5}
//: {6}(378,198)(408,198){7}
//: {8}(412,198)(438,198){9}
//: {10}(442,198)(475,198)(475,235){11}
//: {12}(440,200)(440,210)(441,210)(441,236){13}
//: {14}(410,200)(410,235){15}
//: {16}(376,200)(376,210)(377,210)(377,235){17}
//: {18}(256,200)(256,210)(254,210)(254,232){19}
//: {20}(222,200)(222,210)(220,210)(220,232){21}
input A;    //: /sn:0 {0}(436,236)(436,136){1}
//: {2}(438,134)(470,134)(470,235){3}
//: {4}(434,134)(406,134){5}
//: {6}(402,134)(370,134){7}
//: {8}(366,134)(282,134){9}
//: {10}(278,134)(215,134){11}
//: {12}(211,134)(103,134){13}
//: {14}(213,136)(213,146)(215,146)(215,232){15}
//: {16}(280,136)(280,146)(284,146)(284,232){17}
//: {18}(368,136)(368,146)(372,146)(372,235){19}
//: {20}(404,136)(404,146)(405,146)(405,235){21}
input AcarreoE;    //: /sn:0 {0}(232,46)(232,110)(246,110){1}
//: {2}(250,110)(288,110){3}
//: {4}(292,110)(378,110){5}
//: {6}(382,110)(414,110){7}
//: {8}(418,110)(444,110){9}
//: {10}(448,110)(480,110)(480,235){11}
//: {12}(446,112)(446,236){13}
//: {14}(416,112)(416,122)(415,122)(415,235){15}
//: {16}(380,112)(380,122)(382,122)(382,235){17}
//: {18}(290,112)(290,122)(289,122)(289,232){19}
//: {20}(248,112)(248,122)(249,122)(249,232){21}
output AcarreoS;    //: /sn:0 {0}(247,433)(247,366)(251,366)(251,351){1}
output Suma;    //: /sn:0 {0}(433,432)(433,359)(428,359)(428,344){1}
wire w14;    //: /sn:0 {0}(425,323)(425,301)(410,301)(410,256){1}
wire w20;    //: /sn:0 {0}(475,256)(475,308)(435,308)(435,323){1}
wire w8;    //: /sn:0 {0}(286,253)(286,320)(256,320)(256,330){1}
wire w17;    //: /sn:0 {0}(430,323)(430,300)(441,300)(441,257){1}
wire w2;    //: /sn:0 {0}(217,253)(217,321)(246,321)(246,330){1}
wire w11;    //: /sn:0 {0}(377,256)(377,308)(420,308)(420,323){1}
wire w5;    //: /sn:0 {0}(251,253)(251,330){1}
//: enddecls

  _GGAND3 #(8) g4 (.I0(!AcarreoE), .I1(B), .I2(!A), .Z(w14));   //: @(410,246) /sn:0 /R:3 /w:[ 15 15 21 1 ]
  _GGOR4 #(10) g8 (.I0(w20), .I1(w17), .I2(w14), .I3(w11), .Z(Suma));   //: @(428,334) /sn:0 /R:3 /w:[ 1 0 0 1 1 ]
  _GGAND3 #(8) g3 (.I0(AcarreoE), .I1(!B), .I2(!A), .Z(w11));   //: @(377,246) /sn:0 /R:3 /w:[ 17 17 19 0 ]
  //: IN g13 (AcarreoE) @(232,44) /sn:0 /R:3 /w:[ 0 ]
  _GGAND2 #(6) g2 (.I0(AcarreoE), .I1(A), .Z(w8));   //: @(286,243) /sn:0 /R:3 /w:[ 19 17 0 ]
  _GGAND2 #(6) g1 (.I0(B), .I1(AcarreoE), .Z(w5));   //: @(251,243) /sn:0 /R:3 /w:[ 19 21 0 ]
  //: IN g11 (B) @(96,198) /sn:0 /w:[ 0 ]
  //: joint g16 (AcarreoE) @(248, 110) /w:[ 2 -1 1 20 ]
  //: OUT g10 (Suma) @(433,429) /sn:0 /R:3 /w:[ 0 ]
  //: joint g28 (AcarreoE) @(446, 110) /w:[ 10 -1 9 12 ]
  //: joint g19 (AcarreoE) @(290, 110) /w:[ 4 -1 3 18 ]
  //: joint g27 (B) @(440, 198) /w:[ 10 -1 9 12 ]
  _GGAND3 #(8) g6 (.I0(AcarreoE), .I1(B), .I2(A), .Z(w20));   //: @(475,246) /sn:0 /R:3 /w:[ 11 11 3 0 ]
  _GGOR3 #(8) g7 (.I0(w8), .I1(w5), .I2(w2), .Z(AcarreoS));   //: @(251,341) /sn:0 /R:3 /w:[ 1 1 1 1 ]
  //: OUT g9 (AcarreoS) @(247,430) /sn:0 /R:3 /w:[ 0 ]
  //: joint g15 (B) @(222, 198) /w:[ 2 -1 1 20 ]
  //: joint g20 (A) @(368, 134) /w:[ 7 -1 8 18 ]
  //: joint g17 (B) @(256, 198) /w:[ 4 -1 3 18 ]
  //: joint g25 (B) @(410, 198) /w:[ 8 -1 7 14 ]
  _GGAND3 #(8) g5 (.I0(!AcarreoE), .I1(!B), .I2(A), .Z(w17));   //: @(441,247) /sn:0 /R:3 /w:[ 13 13 0 1 ]
  //: joint g14 (A) @(213, 134) /w:[ 11 -1 12 14 ]
  //: joint g21 (B) @(376, 198) /w:[ 6 -1 5 16 ]
  //: joint g24 (AcarreoE) @(416, 110) /w:[ 8 -1 7 14 ]
  //: joint g23 (A) @(404, 134) /w:[ 5 -1 6 20 ]
  _GGAND2 #(6) g0 (.I0(B), .I1(A), .Z(w2));   //: @(217,243) /sn:0 /R:3 /w:[ 21 15 0 ]
  //: joint g22 (AcarreoE) @(380, 110) /w:[ 6 -1 5 16 ]
  //: joint g26 (A) @(436, 134) /w:[ 2 -1 4 1 ]
  //: IN g12 (A) @(101,134) /sn:0 /w:[ 13 ]
  //: joint g18 (A) @(280, 134) /w:[ 9 -1 10 16 ]

endmodule
//: /netlistEnd

