//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "ETC.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [31:0] w11;    //: /sn:0 {0}(#:149,329)(175,329)(175,297)(210,297){1}
//: {2}(214,297)(347,297){3}
//: {4}(351,297)(#:453,297){5}
//: {6}(349,299)(349,340)(405,340)(405,374){7}
//: {8}(212,299)(212,372){9}
//: {10}(210,374)(192,374)(192,373)(190,373){11}
//: {12}(212,376)(212,408)(130,408)(130,433){13}
reg [2:0] w12;    //: /sn:0 {0}(#:515,66)(515,125){1}
//: {2}(517,127)(577,127){3}
//: {4}(581,127)(602,127)(602,91)(626,91){5}
//: {6}(579,125)(579,52)(625,52){7}
//: {8}(515,129)(#:515,253){9}
reg [31:0] w10;    //: /sn:0 {0}(#:152,241)(175,241)(175,273)(208,273){1}
//: {2}(212,273)(346,273){3}
//: {4}(350,273)(#:453,273){5}
//: {6}(348,271)(#:348,247)(393,247)(393,200){7}
//: {8}(210,271)(210,167){9}
//: {10}(210,163)(210,141)(112,141)(112,122){11}
//: {12}(208,165)(178,165){13}
supply0 w48;    //: /sn:0 {0}(1389,90)(1389,43)(1407,43){1}
//: {2}(1411,43)(1431,43){3}
//: {4}(1435,43)(1547,43){5}
//: {6}(1433,45)(1433,50)(1455,50){7}
//: {8}(1459,50)(1469,50)(1469,53)(1547,53){9}
//: {10}(1457,48)(1457,35){11}
//: {12}(1459,33)(1547,33){13}
//: {14}(1457,31)(1457,15){15}
//: {16}(1459,13)(1547,13){17}
//: {18}(1457,11)(1457,-6){19}
//: {20}(1459,-8)(1469,-8)(1469,-7)(1547,-7){21}
//: {22}(1457,-10)(1457,-29){23}
//: {24}(1459,-31)(1469,-31)(1469,-27)(1547,-27){25}
//: {26}(1457,-33)(1457,-46){27}
//: {28}(1459,-48)(1469,-48)(1469,-47)(1547,-47){29}
//: {30}(1457,-50)(1457,-64){31}
//: {32}(1459,-66)(1469,-66)(1469,-67)(1547,-67){33}
//: {34}(1457,-68)(1457,-83){35}
//: {36}(1459,-85)(1469,-85)(1469,-87)(1547,-87){37}
//: {38}(1457,-87)(1457,-109){39}
//: {40}(1459,-111)(1469,-111)(1469,-107)(1547,-107){41}
//: {42}(1457,-113)(1457,-126){43}
//: {44}(1459,-128)(1469,-128)(1469,-127)(1547,-127){45}
//: {46}(1457,-130)(1457,-152){47}
//: {48}(1459,-154)(1469,-154)(1469,-157)(1547,-157){49}
//: {50}(1457,-156)(1457,-167)(1547,-167){51}
//: {52}(1455,-154)(1445,-154)(1445,-147)(1547,-147){53}
//: {54}(1459,-128)(1449,-128)(1449,-137)(1547,-137){55}
//: {56}(1455,-111)(1445,-111)(1445,-117)(1547,-117){57}
//: {58}(1459,-85)(1449,-85)(1449,-97)(1547,-97){59}
//: {60}(1459,-66)(1449,-66)(1449,-77)(1547,-77){61}
//: {62}(1455,-48)(1445,-48)(1445,-57)(1547,-57){63}
//: {64}(1455,-31)(1445,-31)(1445,-37)(1547,-37){65}
//: {66}(1455,-8)(1445,-8)(1445,-17)(1547,-17){67}
//: {68}(1459,13)(1449,13)(1449,3)(1547,3){69}
//: {70}(1459,33)(1449,33)(1449,23)(1547,23){71}
//: {72}(1457,52)(1457,68){73}
//: {74}(1459,70)(1469,70)(1469,73)(1547,73){75}
//: {76}(1459,70)(1449,70)(1449,63)(1547,63){77}
//: {78}(1457,72)(1457,93){79}
//: {80}(1459,95)(1469,95)(1469,93)(1547,93){81}
//: {82}(1459,95)(1449,95)(1449,83)(1547,83){83}
//: {84}(1457,97)(1457,110){85}
//: {86}(1459,112)(1469,112)(1469,113)(1547,113){87}
//: {88}(1459,112)(1449,112)(1449,103)(1547,103){89}
//: {90}(1457,114)(1457,131){91}
//: {92}(1459,133)(1547,133){93}
//: {94}(1459,133)(1449,133)(1449,123)(1547,123){95}
//: {96}(1457,135)(1457,178){97}
//: {98}(1409,45)(1409,90){99}
supply1 w47;    //: /sn:0 {0}(1313,31)(1313,59)(1397,59){1}
//: {2}(1401,59)(1435,59)(1435,143)(1547,143){3}
//: {4}(1399,61)(1399,90){5}
wire [31:0] w6;    //: /sn:0 {0}(966,307)(1220,307)(1220,344)(1506,344)(#:1506,252)(#:1468,252){1}
wire w7;    //: /sn:0 {0}(1581,279)(1581,288)(1468,288){1}
wire w4;    //: /sn:0 {0}(700,343)(700,353)(666,353)(666,303)(584,303){1}
wire [2:0] w0;    //: /sn:0 {0}(#:1399,96)(#:1399,238){1}
wire w3;    //: /sn:0 {0}(584,285)(684,285)(684,318)(699,318)(699,308){1}
wire [31:0] w1;    //: /sn:0 {0}(#:1553,-12)(1633,-12)(1633,212)(1283,212)(1283,282)(#:1337,282){1}
wire w8;    //: /sn:0 {0}(1564,262)(1564,270)(1468,270){1}
wire [31:0] w2;    //: /sn:0 {0}(#:1069,258)(#:1337,258){1}
wire [31:0] w5;    //: /sn:0 {0}(#:584,267)(676,267)(676,254){1}
//: {2}(678,252)(709,252)(709,241)(739,241){3}
//: {4}(676,250)(676,206)(715,206){5}
//: {6}(674,252)(655,252)(655,258)(1053,258){7}
//: enddecls

  //: comment g61 @(328,146) /sn:0
  //: /line:"Entrada A"
  //: /end
  //: LED g4 (w12) @(632,52) /sn:0 /R:3 /w:[ 7 ] /type:3
  //: DIP g8 (w11) @(111,329) /sn:0 /R:1 /w:[ 0 ] /st:34148 /dn:1
  //: comment g58 @(1336,306) /sn:0
  //: /line:"Esta ALU es para pasr"
  //: /line:"mostrar el negativo en C2"
  //: /end
  //: LED g55 (w8) @(1564,255) /sn:0 /w:[ 0 ] /type:0
  //: joint g51 (w48) @(1457, -128) /w:[ 44 46 54 43 ]
  //: joint g37 (w48) @(1457, 112) /w:[ 86 85 88 90 ]
  //: VDD g34 (w47) @(1324,31) /sn:0 /w:[ 0 ]
  //: LED g3 (w5) @(722,206) /sn:0 /R:3 /w:[ 5 ] /type:3
  //: joint g13 (w10) @(210, 273) /w:[ 2 8 1 -1 ]
  //: LED g2 (w4) @(700,336) /sn:0 /w:[ 0 ] /type:0
  //: comment g59 @(1559,-45) /sn:0
  //: /line:"1 en 32 bits"
  //: /end
  //: LED g1 (w3) @(699,301) /sn:0 /w:[ 1 ] /type:0
  //: LED g11 (w11) @(405,381) /sn:0 /R:2 /w:[ 7 ] /type:3
  //: joint g16 (w11) @(212, 297) /w:[ 2 -1 1 8 ]
  //: joint g50 (w48) @(1457, -111) /w:[ 40 42 56 39 ]
  //: LED g10 (w11) @(130,440) /sn:0 /R:2 /w:[ 13 ] /type:2
  //: joint g28 (w10) @(210, 165) /w:[ -1 10 12 9 ]
  assign w0 = {w48, w47, w48}; //: CONCAT g32  @(1399,95) /sn:0 /R:3 /w:[ 0 0 5 99 ] /dr:1 /tp:0 /drp:1
  //: comment g19 @(664,35) /sn:0
  //: /line:"0 -> AND"
  //: /line:"1 -> OR"
  //: /line:"2 -> Suma"
  //: /line:"6 -> Resta"
  //: /line:"7 -> Compara"
  //: /end
  //: joint g27 (w5) @(676, 252) /w:[ 2 4 6 1 ]
  //: joint g38 (w48) @(1457, 95) /w:[ 80 79 82 84 ]
  //: LED g6 (w10) @(393,193) /sn:0 /w:[ 7 ] /type:3
  //: comment g57 @(789,274) /sn:0
  //: /line:"Salida negativa"
  //: /end
  //: joint g53 (w48) @(1409, 43) /w:[ 2 -1 1 98 ]
  //: DIP g7 (w10) @(114,241) /sn:0 /R:1 /w:[ 0 ] /st:17429 /dn:1
  //: DIP g9 (w12) @(515,56) /sn:0 /w:[ 0 ] /st:2 /dn:1
  _GGNBUF32 #(2) g31 (.I(w5), .Z(w2));   //: @(1059,258) /sn:0 /w:[ 7 0 ]
  //: joint g15 (w11) @(349, 297) /w:[ 4 -1 3 6 ]
  //: comment g20 @(792,171) /sn:0
  //: /line:"Salida"
  //: /end
  //: joint g39 (w47) @(1399, 59) /w:[ 2 -1 1 4 ]
  //: joint g48 (w48) @(1457, -66) /w:[ 32 34 60 31 ]
  //: joint g43 (w48) @(1457, 13) /w:[ 16 18 68 15 ]
  //: comment g62 @(344,417) /sn:0
  //: /line:"Entrada B"
  //: /end
  //: comment g17 @(715,301) /sn:0
  //: /line:"Cero"
  //: /end
  //: LED g25 (w5) @(746,241) /sn:0 /R:3 /w:[ 3 ] /type:1
  //: joint g29 (w11) @(212, 374) /w:[ -1 9 10 12 ]
  //: joint g52 (w48) @(1433, 43) /w:[ 4 -1 3 6 ]
  //: joint g42 (w48) @(1457, 33) /w:[ 12 14 70 11 ]
  //: comment g63 @(3,505) /sn:0
  //: /line:"Gonzalo Caparr�s L�iz"
  //: /end
  //: LED g56 (w7) @(1581,272) /sn:0 /w:[ 0 ] /type:0
  //: LED g5 (w10) @(112,115) /sn:0 /w:[ 11 ] /type:2
  //: joint g14 (w10) @(348, 273) /w:[ 4 6 3 -1 ]
  //: joint g47 (w48) @(1457, -48) /w:[ 28 30 62 27 ]
  //: joint g44 (w48) @(1457, -8) /w:[ 20 22 66 19 ]
  //: joint g36 (w48) @(1457, 133) /w:[ 92 91 94 96 ]
  //: comment g21 @(490,15) /sn:0
  //: /line:"Control"
  //: /end
  //: LED g24 (w12) @(633,91) /sn:0 /R:3 /w:[ 5 ] /type:1
  //: joint g41 (w48) @(1457, 50) /w:[ 8 10 7 72 ]
  //: LED g23 (w11) @(183,373) /sn:0 /R:1 /w:[ 11 ] /type:1
  //: comment g60 @(1275,69) /sn:0
  //: /line:"Senal de control"
  //: /line:"para sumar"
  //: /end
  //: LED g54 (w6) @(959,307) /sn:0 /R:1 /w:[ 0 ] /type:3
  //: joint g40 (w48) @(1457, 70) /w:[ 74 73 76 78 ]
  //: joint g46 (w48) @(1457, -31) /w:[ 24 26 64 23 ]
  //: joint g45 (w48) @(1457, -154) /w:[ 48 50 52 47 ]
  //: GROUND g35 (w48) @(1457,184) /sn:0 /w:[ 97 ]
  ALU g0 (.C(w12), .B(w11), .A(w10), .Sa(w5), .Overflow(w4), .Cero(w3));   //: @(454, 254) /sz:(129, 64) /sn:0 /p:[ Ti0>9 Li0>5 Li1>5 Ro0<0 Ro1<1 Ro2<0 ]
  //: LED g22 (w10) @(171,165) /sn:0 /R:1 /w:[ 13 ] /type:1
  //: joint g26 (w12) @(579, 127) /w:[ 4 6 3 -1 ]
  //: joint g12 (w12) @(515, 127) /w:[ 2 1 -1 8 ]
  //: comment g18 @(718,338) /sn:0
  //: /line:"Overflow"
  //: /end
  assign w1 = {w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w48, w47}; //: CONCAT g33  @(1552,-12) /sn:0 /w:[ 0 51 49 53 55 45 57 41 59 37 61 33 63 29 65 25 67 21 69 17 71 13 5 9 77 75 83 81 89 87 95 93 3 ] /dr:0 /tp:0 /drp:1
  ALU g30 (.C(w0), .A(w2), .B(w1), .Cero(w8), .Overflow(w7), .Sa(w6));   //: @(1338, 239) /sz:(129, 64) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Ro0<1 Ro1<1 Ro2<1 ]
  //: joint g49 (w48) @(1457, -85) /w:[ 36 38 58 35 ]

endmodule
//: /netlistEnd

//: /netlistBegin FlipFlopD
module FlipFlopD(Reloj, nQ, Q, D, W);
//: interface  /sz:(129, 78) /bd:[ Li0>Reloj(51/78) Li1>D(25/78) Bi0>W(71/129) Ro0<nQ(54/78) Ro1<Q(27/78) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output Q;    //: /sn:0 {0}(458,116)(551,116)(551,109)(566,109){1}
output nQ;    //: /sn:0 {0}(458,135)(536,135)(536,191)(551,191){1}
input D;    //: /sn:0 {0}(47,98)(158,98)(158,110)(188,110){1}
input Reloj;    //: /sn:0 {0}(46,293)(81,293)(81,281)(96,281){1}
input W;    //: /sn:0 {0}(374,327)(374,265){1}
//: {2}(374,261)(374,237)(359,237)(359,224){3}
//: {4}(372,263)(169,263)(169,224){5}
wire w0;    //: /sn:0 {0}(112,281)(139,281)(139,293)(162,293){1}
//: {2}(166,293)(196,293)(196,281)(207,281){3}
//: {4}(164,291)(164,224){5}
wire w3;    //: /sn:0 {0}(280,127)(265,127){1}
wire w1;    //: /sn:0 {0}(167,203)(167,125)(188,125){1}
wire w2;    //: /sn:0 {0}(265,108)(362,108)(362,118)(381,118){1}
wire w5;    //: /sn:0 {0}(357,203)(357,133)(381,133){1}
wire w9;    //: /sn:0 {0}(354,224)(354,281)(223,281){1}
//: enddecls

  _GGAND2 #(6) g4 (.I0(w0), .I1(W), .Z(w1));   //: @(167,213) /sn:0 /R:1 /w:[ 5 5 0 ]
  //: IN g8 (Reloj) @(44,293) /sn:0 /w:[ 0 ]
  //: joint g13 (w0) @(164, 293) /w:[ 2 4 1 -1 ]
  //: OUT g3 (nQ) @(548,191) /sn:0 /w:[ 1 ]
  //: OUT g2 (Q) @(563,109) /sn:0 /w:[ 1 ]
  LatchD g1 (.C(w5), .D(w2), .nQ(nQ), .Q(Q));   //: @(382, 104) /sz:(75, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  //: joint g11 (W) @(374, 263) /w:[ -1 2 4 1 ]
  _GGNBUF #(2) g10 (.I(Reloj), .Z(w0));   //: @(102,281) /sn:0 /w:[ 1 0 ]
  _GGNBUF #(2) g6 (.I(w0), .Z(w9));   //: @(213,281) /sn:0 /w:[ 3 1 ]
  //: IN g7 (D) @(45,98) /sn:0 /w:[ 0 ]
  //: IN g9 (W) @(374,329) /sn:0 /R:1 /w:[ 0 ]
  _GGAND2 #(6) g5 (.I0(w9), .I1(W), .Z(w5));   //: @(357,213) /sn:0 /R:1 /w:[ 0 3 0 ]
  LatchD g0 (.C(w1), .D(D), .nQ(w3), .Q(w2));   //: @(189, 96) /sz:(75, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  //: comment g12 @(343,29) /sn:0
  //: /line:"Flanco ascendente"
  //: /end

endmodule
//: /netlistEnd

//: /netlistBegin LatchSR
module LatchSR(C, Q, S, R, nQ);
//: interface  /sz:(81, 64) /bd:[ Li0>S(11/64) Li1>R(46/64) Li2>C(28/64) Ro0<Q(20/64) Ro1<nQ(40/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output nQ;    //: /sn:0 {0}(435,245)(500,245){1}
//: {2}(504,245)(561,245){3}
//: {4}(502,243)(502,137)(412,137)(412,122)(422,122){5}
output Q;    //: /sn:0 {0}(443,120)(505,120)(505,112)(521,112){1}
//: {2}(525,112)(563,112){3}
//: {4}(523,114)(523,227)(404,227)(404,242)(414,242){5}
input R;    //: /sn:0 {0}(156,97)(304,97)(304,114)(319,114){1}
input C;    //: /sn:0 {0}(173,192)(258,192){1}
//: {2}(260,190)(260,119)(319,119){3}
//: {4}(260,194)(260,258)(307,258){5}
input S;    //: /sn:0 {0}(196,295)(292,295)(292,263)(307,263){1}
wire w2;    //: /sn:0 {0}(340,117)(422,117){1}
wire w5;    //: /sn:0 {0}(328,261)(399,261)(399,247)(414,247){1}
//: enddecls

  //: IN g8 (C) @(171,192) /sn:0 /w:[ 0 ]
  //: OUT g4 (Q) @(560,112) /sn:0 /w:[ 3 ]
  _GGNOR2 #(4) g3 (.I0(Q), .I1(w5), .Z(nQ));   //: @(425,245) /sn:0 /w:[ 5 1 0 ]
  _GGNOR2 #(4) g2 (.I0(w2), .I1(nQ), .Z(Q));   //: @(433,120) /sn:0 /w:[ 1 5 0 ]
  _GGAND2 #(6) g1 (.I0(C), .I1(S), .Z(w5));   //: @(318,261) /sn:0 /w:[ 5 1 0 ]
  //: joint g11 (Q) @(523, 112) /w:[ 2 -1 1 4 ]
  //: joint g10 (nQ) @(502, 245) /w:[ 2 4 1 -1 ]
  //: IN g6 (S) @(194,295) /sn:0 /w:[ 0 ]
  //: joint g9 (C) @(260, 192) /w:[ -1 2 1 4 ]
  //: IN g7 (R) @(154,97) /sn:0 /w:[ 0 ]
  //: OUT g5 (nQ) @(558,245) /sn:0 /w:[ 3 ]
  _GGAND2 #(6) g0 (.I0(R), .I1(C), .Z(w2));   //: @(330,117) /sn:0 /w:[ 1 3 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FlipFlopT
module FlipFlopT(Q, nQ, Reloj, T);
//: interface  /sz:(106, 65) /bd:[ Li0>T(25/65) Li1>Reloj(45/65) Ro0<Q(17/65) Ro1<nQ(37/65) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output nQ;    //: /sn:0 {0}(172,254)(162,254)(162,284)(385,284)(385,234){1}
//: {2}(387,232)(436,232)(436,236)(447,236){3}
//: {4}(383,232)(374,232)(374,231)(368,231){5}
//: {6}(366,229)(366,163)(301,163)(301,149)(313,149){7}
//: {8}(364,231)(346,231)(346,232)(331,232){9}
output Q;    //: /sn:0 {0}(334,147)(365,147)(365,148)(391,148){1}
//: {2}(395,148)(445,148){3}
//: {4}(393,146)(393,93)(179,93)(179,117)(183,117){5}
//: {6}(393,150)(393,215)(306,215)(306,229)(310,229){7}
input T;    //: /sn:0 {0}(41,125)(98,125){1}
//: {2}(102,125)(147,125)(147,122)(183,122){3}
//: {4}(100,127)(100,249)(172,249){5}
input Reloj;    //: /sn:0 {0}(57,174)(141,174)(141,178)(155,178){1}
//: {2}(157,176)(157,127)(183,127){3}
//: {4}(157,180)(157,244)(172,244){5}
wire w6;    //: /sn:0 {0}(193,249)(295,249)(295,234)(310,234){1}
wire w2;    //: /sn:0 {0}(204,122)(298,122)(298,144)(313,144){1}
//: enddecls

  _GGNOR2 #(4) g8 (.I0(Q), .I1(w6), .Z(nQ));   //: @(321,232) /sn:0 /w:[ 7 1 9 ]
  //: OUT g4 (Q) @(442,148) /sn:0 /w:[ 3 ]
  //: OUT g3 (nQ) @(444,236) /sn:0 /w:[ 3 ]
  //: comment g13 @(179,46) /sn:0
  //: /line:"Como pone en internet(no funciona)"
  //: /end
  //: joint g2 (T) @(100, 125) /w:[ 2 -1 1 4 ]
  //: IN g1 (Reloj) @(55,174) /sn:0 /w:[ 0 ]
  //: joint g11 (nQ) @(366, 231) /w:[ 5 6 8 -1 ]
  //: joint g10 (Q) @(393, 148) /w:[ 2 4 1 6 ]
  _GGAND3 #(8) g6 (.I0(Reloj), .I1(T), .I2(nQ), .Z(w6));   //: @(183,249) /sn:0 /w:[ 5 5 0 0 ]
  //: joint g9 (Reloj) @(157, 178) /w:[ -1 2 1 4 ]
  _GGNOR2 #(4) g7 (.I0(w2), .I1(nQ), .Z(Q));   //: @(324,147) /sn:0 /w:[ 1 7 0 ]
  _GGAND3 #(8) g5 (.I0(Q), .I1(T), .I2(Reloj), .Z(w2));   //: @(194,122) /sn:0 /w:[ 5 3 3 0 ]
  //: IN g0 (T) @(39,125) /sn:0 /w:[ 0 ]
  //: joint g12 (nQ) @(385, 232) /w:[ 2 -1 4 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin FlipFlopSR
module FlipFlopSR(nQ, R, S, Reloj, Q);
//: interface  /sz:(134, 64) /bd:[ Li0>S(14/64) Li1>Reloj(32/64) Li2>R(52/64) Ro0<Q(27/64) Ro1<nQ(44/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output nQ;    //: /sn:0 {0}(453,123)(550,123)(550,157)(565,157){1}
output Q;    //: /sn:0 {0}(453,103)(545,103)(545,100)(560,100){1}
input R;    //: /sn:0 {0}(58,157)(154,157)(154,130)(179,130){1}
input Reloj;    //: /sn:0 {0}(56,266)(89,266)(89,238)(104,238){1}
input S;    //: /sn:0 {0}(56,92)(131,92)(131,95)(179,95){1}
wire w7;    //: /sn:0 {0}(287,255)(355,255)(355,111)(370,111){1}
wire w4;    //: /sn:0 {0}(262,104)(273,104)(273,94)(370,94){1}
wire w0;    //: /sn:0 {0}(179,112)(148,112)(148,264){1}
//: {2}(150,266)(160,266)(160,255)(271,255){3}
//: {4}(146,266)(128,266)(128,238)(120,238){5}
wire w3;    //: /sn:0 {0}(262,124)(331,124)(331,129)(370,129){1}
//: enddecls

  //: OUT g8 (nQ) @(562,157) /sn:0 /w:[ 1 ]
  _GGNBUF #(2) g4 (.I(Reloj), .Z(w0));   //: @(110,238) /sn:0 /w:[ 1 5 ]
  //: IN g3 (R) @(56,157) /sn:0 /w:[ 0 ]
  //: IN g2 (S) @(54,92) /sn:0 /w:[ 0 ]
  LatchSR g1 (.C(w7), .R(w3), .S(w4), .nQ(nQ), .Q(Q));   //: @(371, 83) /sz:(81, 64) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Ro0<0 Ro1<0 ]
  //: comment g10 @(266,23) /sn:0
  //: /line:"Flancao ascendente"
  //: /end
  //: IN g6 (Reloj) @(54,266) /sn:0 /w:[ 0 ]
  //: joint g9 (w0) @(148, 266) /w:[ 2 1 4 -1 ]
  //: OUT g7 (Q) @(557,100) /sn:0 /w:[ 1 ]
  _GGNBUF #(2) g5 (.I(w0), .Z(w7));   //: @(277,255) /sn:0 /w:[ 3 0 ]
  LatchSR g0 (.C(w0), .R(R), .S(S), .nQ(w3), .Q(w4));   //: @(180, 84) /sz:(81, 64) /sn:0 /p:[ Li0>0 Li1>1 Li2>1 Ro0<0 Ro1<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin ALU
module ALU(Sa, Cero, B, A, C, Overflow);
//: interface  /sz:(129, 64) /bd:[ Ti0>C[2:0](61/129) Li0>B[31:0](43/64) Li1>A[31:0](19/64) Ro0<Sa[31:0](13/64) Ro1<Overflow(49/64) Ro2<Cero(31/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [31:0] A;    //: /sn:0 {0}(#:-133,-78)(-114,-78)(-114,-226)(#:71,-226){1}
supply0 w54;    //: /sn:0 {0}(476,-314)(476,-361){1}
//: {2}(478,-363)(509,-363){3}
//: {4}(476,-365)(476,-372)(509,-372){5}
//: {6}(478,-363)(468,-363)(468,-353)(509,-353){7}
output Cero;    //: /sn:0 {0}(1741,915)(1731,915)(1731,916)(1675,916){1}
output Overflow;    //: /sn:0 {0}(383,2652)(383,2708)(413,2708){1}
output [31:0] Sa;    //: /sn:0 {0}(#:1263,925)(1138,925)(1138,1133){1}
//: {2}(1140,1135)(1325,1135){3}
//: {4}(1136,1135)(#:1034,1135){5}
input [2:0] C;    //: /sn:0 {0}(#:537,2331)(537,2253){1}
//: {2}(539,2251)(716,2251)(716,2169){3}
//: {4}(716,2165)(716,2079){5}
//: {6}(716,2075)(716,1998){7}
//: {8}(716,1994)(716,1913){9}
//: {10}(716,1909)(716,1828){11}
//: {12}(716,1824)(716,1748){13}
//: {14}(716,1744)(716,1661){15}
//: {16}(716,1657)(716,1575){17}
//: {18}(716,1571)(716,1489){19}
//: {20}(716,1485)(716,1416){21}
//: {22}(716,1412)(716,1340){23}
//: {24}(716,1336)(716,1238){25}
//: {26}(716,1234)(716,1151){27}
//: {28}(716,1147)(716,1094){29}
//: {30}(716,1090)(716,992){31}
//: {32}(716,988)(716,898){33}
//: {34}(716,894)(716,826){35}
//: {36}(716,822)(716,741){37}
//: {38}(716,737)(716,657){39}
//: {40}(716,653)(716,561){41}
//: {42}(716,557)(716,461){43}
//: {44}(716,457)(716,373){45}
//: {46}(716,369)(716,284){47}
//: {48}(716,280)(716,197){49}
//: {50}(716,193)(716,140)(717,140)(717,106){51}
//: {52}(717,102)(717,6){53}
//: {54}(717,2)(717,-80){55}
//: {56}(717,-84)(717,-172){57}
//: {58}(717,-176)(717,-277){59}
//: {60}(717,-281)(717,-536)(575,-536){61}
//: {62}(573,-538)(573,-543)(541,-543)(#:541,-546){63}
//: {64}(573,-534)(573,-526)(541,-526)(#:541,-515){65}
//: {66}(715,-279)(431,-279)(431,-257){67}
//: {68}(715,-174)(432,-174)(432,-160){69}
//: {70}(715,-82)(433,-82)(433,-63){71}
//: {72}(715,4)(434,4)(#:434,27){73}
//: {74}(715,104)(435,104)(#:435,118){75}
//: {76}(714,195)(436,195)(#:436,211){77}
//: {78}(714,282)(437,282)(#:437,299){79}
//: {80}(714,371)(438,371)(#:438,393){81}
//: {82}(714,459)(439,459)(#:439,481){83}
//: {84}(714,559)(442,559)(#:442,572){85}
//: {86}(714,655)(509,655)(509,645)(452,645)(#:452,661){87}
//: {88}(714,739)(462,739)(#:462,744){89}
//: {90}(714,824)(444,824)(#:444,829){91}
//: {92}(714,896)(440,896)(#:440,913){93}
//: {94}(714,990)(436,990)(#:436,999){95}
//: {96}(714,1092)(521,1092)(521,1070)(444,1070)(#:444,1082){97}
//: {98}(714,1149)(439,1149)(#:439,1170){99}
//: {100}(714,1236)(459,1236)(#:459,1263){101}
//: {102}(714,1338)(515,1338)(515,1329)(471,1329)(#:471,1343){103}
//: {104}(714,1414)(454,1414)(#:454,1424){105}
//: {106}(714,1487)(451,1487)(#:451,1507){107}
//: {108}(714,1573)(444,1573)(#:444,1592){109}
//: {110}(714,1659)(439,1659)(#:439,1673){111}
//: {112}(714,1746)(451,1746)(#:451,1753){113}
//: {114}(714,1826)(444,1826)(#:444,1839){115}
//: {116}(714,1911)(442,1911)(#:442,1920){117}
//: {118}(714,1996)(429,1996)(#:429,2005){119}
//: {120}(714,2077)(454,2077)(#:454,2093){121}
//: {122}(714,2167)(440,2167)(#:440,2172){123}
//: {124}(535,2251)(461,2251)(#:461,2256){125}
input [31:0] B;    //: /sn:0 {0}(#:-653,763)(#:-290,763){1}
supply0 w49;    //: /sn:0 {0}(467,2432)(441,2432){1}
//: {2}(439,2430)(439,2423)(467,2423){3}
//: {4}(439,2434)(439,2446)(449,2446){5}
//: {6}(451,2444)(451,2442)(467,2442){7}
//: {8}(451,2448)(451,2461){9}
//: {10}(453,2463)(467,2463){11}
//: {12}(451,2465)(451,2498){13}
wire w32;    //: /sn:0 {0}(332,2481)(297,2481){1}
//: {2}(293,2481)(98,2481)(98,2409){3}
//: {4}(100,2407)(110,2407)(110,2412)(292,2412){5}
//: {6}(98,2405)(98,2394){7}
//: {8}(100,2392)(110,2392)(110,2395)(292,2395){9}
//: {10}(98,2390)(98,-71)(77,-71){11}
//: {12}(295,2483)(295,2563)(371,2563)(371,2607){13}
wire w45;    //: /sn:0 {0}(-284,728)(355,728)(355,781)(395,781){1}
wire w73;    //: /sn:0 {0}(1028,1050)(981,1050)(981,331)(459,331){1}
wire w96;    //: /sn:0 {0}(1028,1280)(857,1280)(857,2288)(483,2288){1}
wire w214;    //: /sn:0 {0}(384,1544)(304,1544)(304,818)(-284,818){1}
wire w244;    //: /sn:0 {0}(394,2293)(257,2293)(257,908)(-284,908){1}
wire w122;    //: /sn:0 {0}(398,-98)(398,-79)(370,-79)(370,-70)(398,-70)(398,-63){1}
wire w134;    //: /sn:0 {0}(369,248)(275,248)(275,668)(-284,668){1}
wire w166;    //: /sn:0 {0}(377,866)(350,866)(350,738)(-284,738){1}
wire w203;    //: /sn:0 {0}(419,1424)(419,1415)(437,1415)(437,1405){1}
wire w220;    //: /sn:0 {0}(375,1957)(279,1957)(279,868)(-284,868){1}
wire w141;    //: /sn:0 {0}(403,361)(403,378)(394,378)(394,385)(403,385)(403,393){1}
wire w14;    //: /sn:0 {0}(77,-251)(167,-251)(167,851)(377,851){1}
wire w16;    //: /sn:0 {0}(77,-231)(158,-231)(158,1021)(369,1021){1}
wire w56;    //: /sn:0 {0}(372,1710)(294,1710)(294,838)(-284,838){1}
wire w179;    //: /sn:0 {0}(409,1082)(409,1076)(402,1076)(402,1061){1}
wire w4;    //: /sn:0 {0}(77,-351)(214,-351)(214,-41)(366,-41){1}
wire w19;    //: /sn:0 {0}(392,1285)(144,1285)(144,-201)(77,-201){1}
wire w81;    //: /sn:0 {0}(1028,1130)(943,1130)(943,1031)(458,1031){1}
wire w89;    //: /sn:0 {0}(461,1705)(789,1705)(789,1210)(1028,1210){1}
wire w195;    //: /sn:0 {0}(473,1785)(798,1785)(798,1220)(1028,1220){1}
wire w38;    //: /sn:0 {0}(368,155)(265,155)(265,658)(-284,658){1}
wire w152;    //: /sn:0 {0}(371,430)(301,430)(301,688)(-284,688){1}
wire w3;    //: /sn:0 {0}(77,-361)(218,-361)(218,-138)(365,-138){1}
wire w0;    //: /sn:0 {0}(362,-334)(325,-334)(325,-362){1}
//: {2}(327,-364)(347,-364){3}
//: {4}(325,-366)(325,-379){5}
//: {6}(327,-381)(347,-381){7}
//: {8}(323,-381)(77,-381){9}
wire w151;    //: /sn:0 {0}(377,1629)(298,1629)(298,828)(-284,828){1}
wire w128;    //: /sn:0 {0}(1269,1060)(1609,1060)(1609,984)(1654,984){1}
wire w127;    //: /sn:0 {0}(1269,1050)(1599,1050)(1599,979)(1654,979){1}
wire w120;    //: /sn:0 {0}(1028,1000)(1000,1000)(1000,-128)(454,-128){1}
wire w233;    //: /sn:0 {0}(405,2172)(405,2165)(420,2165)(420,2155){1}
wire w240;    //: /sn:0 {0}(1028,1270)(846,1270)(846,2204)(462,2204){1}
wire w133;    //: /sn:0 {0}(-284,708)(320,708)(320,609)(375,609){1}
wire w104;    //: /sn:0 {0}(396,-288)(396,-274)(385,-274)(385,-266)(396,-266)(396,-257){1}
wire w111;    //: /sn:0 {0}(368,-378)(428,-378)(428,-403)(509,-403){1}
wire w168;    //: /sn:0 {0}(1028,1110)(954,1110)(954,861)(466,861){1}
wire w204;    //: /sn:0 {0}(1028,1170)(750,1170)(750,1375)(493,1375){1}
wire w75;    //: /sn:0 {0}(1028,1070)(973,1070)(973,513)(461,513){1}
wire w209;    //: /sn:0 {0}(416,1507)(416,1495)(420,1495)(420,1486){1}
wire w67;    //: /sn:0 {0}(1028,990)(1005,990)(1005,-225)(453,-225){1}
wire w119;    //: /sn:0 {0}(400,118)(400,106)(387,106)(387,97)(400,97)(400,89){1}
wire w90;    //: /sn:0 {0}(1269,910)(1513,910)(1513,909)(1654,909){1}
wire w215;    //: /sn:0 {0}(409,1592)(409,1574)(417,1574)(417,1569){1}
wire w156;    //: /sn:0 {0}(1028,1090)(965,1090)(965,693)(474,693){1}
wire w167;    //: /sn:0 {0}(405,913)(405,904)(396,904)(396,896)(410,896)(410,891){1}
wire w41;    //: /sn:0 {0}(313,2415)(387,2415)(387,2404)(467,2404){1}
wire w36;    //: /sn:0 {0}(366,-26)(252,-26)(252,638)(-284,638){1}
wire w20;    //: /sn:0 {0}(77,-191)(139,-191)(139,1365)(404,1365){1}
wire w23;    //: /sn:0 {0}(377,1614)(129,1614)(129,-161)(77,-161){1}
wire w124;    //: /sn:0 {0}(1028,1020)(992,1020)(992,59)(456,59){1}
wire w174;    //: /sn:0 {0}(1028,1120)(949,1120)(949,945)(462,945){1}
wire w82;    //: /sn:0 {0}(1028,1140)(939,1140)(939,1114)(466,1114){1}
wire w126;    //: /sn:0 {0}(1028,1010)(996,1010)(996,-31)(455,-31){1}
wire w74;    //: /sn:0 {0}(1028,1060)(977,1060)(977,425)(460,425){1}
wire w125;    //: /sn:0 {0}(399,-1)(399,13)(371,13)(371,19)(399,19)(399,27){1}
wire w91;    //: /sn:0 {0}(466,1871)(806,1871)(806,1230)(1028,1230){1}
wire w35;    //: /sn:0 {0}(365,-123)(247,-123)(247,628)(-284,628){1}
wire w8;    //: /sn:0 {0}(77,-311)(195,-311)(195,321)(370,321){1}
wire w103;    //: /sn:0 {0}(551,-509)(551,-467)(552,-467)(552,-411){1}
wire w101;    //: /sn:0 {0}(1269,970)(1542,970)(1542,939)(1654,939){1}
wire w192;    //: /sn:0 {0}(461,1202)(724,1202)(724,1150)(1028,1150){1}
wire w71;    //: /sn:0 {0}(1028,1030)(988,1030)(988,150)(457,150){1}
wire w202;    //: /sn:0 {0}(404,1380)(313,1380)(313,798)(-284,798){1}
wire w238;    //: /sn:0 {0}(373,2209)(261,2209)(261,898)(-284,898){1}
wire w22;    //: /sn:0 {0}(384,1529)(133,1529)(133,-171)(77,-171){1}
wire w17;    //: /sn:0 {0}(377,1104)(153,1104)(153,-221)(77,-221){1}
wire w117;    //: /sn:0 {0}(1269,1010)(1563,1010)(1563,959)(1654,959){1}
wire w53;    //: /sn:0 {0}(387,1461)(308,1461)(308,808)(-284,808){1}
wire w84;    //: /sn:0 {0}(1028,1160)(739,1160)(739,1295)(481,1295){1}
wire w172;    //: /sn:0 {0}(-284,748)(344,748)(344,950)(373,950){1}
wire w211;    //: /sn:0 {0}(407,1920)(407,1908)(410,1908)(410,1901){1}
wire w228;    //: /sn:0 {0}(1028,1250)(823,1250)(823,2037)(451,2037){1}
wire w12;    //: /sn:0 {0}(385,683)(177,683)(177,-271)(77,-271){1}
wire w113;    //: /sn:0 {0}(397,-195)(397,-180)(383,-180)(383,-172)(397,-172)(397,-160){1}
wire w44;    //: /sn:0 {0}(-284,718)(326,718)(326,698)(385,698){1}
wire w2;    //: /sn:0 {0}(396,-350)(396,-462){1}
//: {2}(398,-464)(528,-464){3}
//: {4}(530,-466)(530,-496)(531,-496)(531,-509){5}
//: {6}(530,-462)(530,-411){7}
//: {8}(394,-464)(284,-464)(284,-353)(309,-353)(309,-330){9}
wire w115;    //: /sn:0 {0}(1269,990)(1554,990)(1554,949)(1654,949){1}
wire w83;    //: /sn:0 {0}(1269,870)(1548,870)(1548,889)(1654,889){1}
wire w77;    //: /sn:0 {0}(1269,850)(1569,850)(1569,879)(1654,879){1}
wire w226;    //: /sn:0 {0}(362,2042)(273,2042)(273,878)(-284,878){1}
wire w78;    //: /sn:0 {0}(1028,1100)(960,1100)(960,776)(484,776){1}
wire w10;    //: /sn:0 {0}(372,503)(186,503)(186,-291)(77,-291){1}
wire w27;    //: /sn:0 {0}(375,1942)(114,1942)(114,-121)(77,-121){1}
wire w190;    //: /sn:0 {0}(372,1207)(326,1207)(326,778)(-284,778){1}
wire w95;    //: /sn:0 {0}(1269,940)(1528,940)(1528,924)(1654,924){1}
wire w52;    //: /sn:0 {0}(1028,1290)(869,1290)(869,2426)(521,2426){1}
wire w86;    //: /sn:0 {0}(1028,1180)(762,1180)(762,1456)(476,1456){1}
wire w80;    //: /sn:0 {0}(213,2538)(142,2538){1}
//: {2}(138,2538)(97,2538){3}
//: {4}(93,2538)(-18,2538)(-18,2412){5}
//: {6}(-16,2410)(-6,2410)(-6,2417)(292,2417){7}
//: {8}(-18,2408)(-18,918)(-284,918){9}
//: {10}(-20,2410)(-30,2410)(-30,2400)(292,2400){11}
//: {12}(95,2540)(95,2588)(392,2588)(392,2607){13}
//: {14}(140,2540)(140,2556)(157,2556){15}
wire w29;    //: /sn:0 {0}(387,2115)(107,2115)(107,-101)(77,-101){1}
wire w155;    //: /sn:0 {0}(427,744)(427,735)(418,735)(418,723){1}
wire w178;    //: /sn:0 {0}(369,1036)(338,1036)(338,758)(-284,758){1}
wire w50;    //: /sn:0 {0}(1269,780)(1628,780)(1628,844)(1654,844){1}
wire w147;    //: /sn:0 {0}(407,572)(407,562)(399,562)(399,553)(405,553)(405,543){1}
wire w42;    //: /sn:0 {0}(-284,698)(311,698)(311,518)(372,518){1}
wire w6;    //: /sn:0 {0}(77,-331)(204,-331)(204,140)(368,140){1}
wire w93;    //: /sn:0 {0}(1654,914)(1517,914)(1517,920)(1269,920){1}
wire w7;    //: /sn:0 {0}(77,-321)(199,-321)(199,233)(369,233){1}
wire w99;    //: /sn:0 {0}(1269,960)(1536,960)(1536,934)(1654,934){1}
wire w175;    //: /sn:0 {0}(416,1753)(416,1744)(405,1744)(405,1735){1}
wire w112;    //: /sn:0 {0}(77,-371)(221,-371)(221,-235)(364,-235){1}
wire w61;    //: /sn:0 {0}(387,2130)(267,2130)(267,888)(-284,888){1}
wire w135;    //: /sn:0 {0}(402,299)(402,286)(394,286)(394,279)(402,279)(402,273){1}
wire w15;    //: /sn:0 {0}(373,935)(163,935)(163,-241)(77,-241){1}
wire w216;    //: /sn:0 {0}(473,1539)(771,1539)(771,1190)(1028,1190){1}
wire w69;    //: /sn:0 {0}(1269,820)(1591,820)(1591,864)(1654,864){1}
wire w239;    //: /sn:0 {0}(426,2256)(426,2244)(406,2244)(406,2234){1}
wire w207;    //: /sn:0 {0}(377,1876)(283,1876)(283,858)(-284,858){1}
wire w51;    //: /sn:0 {0}(392,1300)(319,1300)(319,788)(-284,788){1}
wire w109;    //: /sn:0 {0}(364,-220)(242,-220)(242,618)(-284,618){1}
wire w129;    //: /sn:0 {0}(401,211)(401,193)(391,193)(391,185)(401,185)(401,180){1}
wire w114;    //: /sn:0 {0}(1269,980)(1548,980)(1548,944)(1654,944){1}
wire w97;    //: /sn:0 {0}(1269,950)(1532,950)(1532,929)(1654,929){1}
wire w64;    //: /sn:0 {0}(1269,810)(1599,810)(1599,859)(1654,859){1}
wire w66;    //: /sn:0 {0}(563,-369)(1010,-369)(1010,980)(1028,980){1}
wire w37;    //: /sn:0 {0}(367,64)(257,64)(257,648)(-284,648){1}
wire w245;    //: /sn:0 {0}(427,2318)(427,2374)(366,2374)(366,2465){1}
wire w63;    //: /sn:0 {0}(1269,800)(1608,800)(1608,854)(1654,854){1}
wire w34;    //: /sn:0 {0}(537,2337)(537,2365)(499,2365)(499,2384){1}
wire w234;    //: /sn:0 {0}(1028,1260)(834,1260)(834,2125)(476,2125){1}
wire w159;    //: /sn:0 {0}(466,1624)(780,1624)(780,1200)(1028,1200){1}
wire w43;    //: /sn:0 {0}(1269,770)(1639,770)(1639,839)(1654,839){1}
wire w87;    //: /sn:0 {0}(1269,890)(1532,890)(1532,899)(1654,899){1}
wire w157;    //: /sn:0 {0}(404,1673)(404,1662)(410,1662)(410,1654){1}
wire w102;    //: /sn:0 {0}(541,-509)(541,-411){1}
wire w76;    //: /sn:0 {0}(1028,1080)(969,1080)(969,604)(464,604){1}
wire w21;    //: /sn:0 {0}(77,-181)(136,-181)(136,1446)(387,1446){1}
wire w100;    //: /sn:0 {0}(431,-321)(455,-321)(455,-340){1}
//: {2}(457,-342)(509,-342){3}
//: {4}(455,-344)(455,-383)(509,-383){5}
wire w31;    //: /sn:0 {0}(394,2278)(101,2278)(101,-81)(77,-81){1}
wire w130;    //: /sn:0 {0}(1269,1070)(1625,1070)(1625,989)(1654,989){1}
wire w28;    //: /sn:0 {0}(362,2027)(111,2027)(111,-111)(77,-111){1}
wire w24;    //: /sn:0 {0}(77,-151)(126,-151)(126,1695)(372,1695){1}
wire w1;    //: /sn:0 {0}(547,2337)(547,2371)(510,2371)(510,2384){1}
wire w161;    //: /sn:0 {0}(409,829)(409,815)(428,815)(428,806){1}
wire w184;    //: /sn:0 {0}(377,1119)(332,1119)(332,768)(-284,768){1}
wire w221;    //: /sn:0 {0}(394,2005)(394,1989)(408,1989)(408,1982){1}
wire w140;    //: /sn:0 {0}(370,336)(289,336)(289,678)(-284,678){1}
wire w25;    //: /sn:0 {0}(77,-141)(123,-141)(123,1775)(384,1775){1}
wire w116;    //: /sn:0 {0}(1269,1000)(1559,1000)(1559,954)(1654,954){1}
wire w227;    //: /sn:0 {0}(419,2093)(419,2079)(395,2079)(395,2067){1}
wire w65;    //: /sn:0 {0}(467,2453)(448,2453){1}
//: {2}(444,2453)(426,2453){3}
//: {4}(424,2451)(424,2412)(467,2412){5}
//: {6}(424,2455)(424,2492){7}
//: {8}(422,2494)(401,2494){9}
//: {10}(424,2496)(424,2558)(414,2558)(414,2607){11}
//: {12}(446,2455)(446,2488)(437,2488)(437,2526)(620,2526)(620,-317)(499,-317)(499,-332)(509,-332){13}
wire w98;    //: /sn:0 {0}(288,-301)(256,-301){1}
wire w121;    //: /sn:0 {0}(1269,1030)(1575,1030)(1575,969)(1654,969){1}
wire w118;    //: /sn:0 {0}(1269,1020)(1568,1020)(1568,964)(1654,964){1}
wire w40;    //: /sn:0 {0}(313,2398)(445,2398)(445,2392)(467,2392){1}
wire w92;    //: /sn:0 {0}(1028,1240)(815,1240)(815,1952)(464,1952){1}
wire w18;    //: /sn:0 {0}(372,1192)(148,1192)(148,-211)(77,-211){1}
wire w68;    //: /sn:0 {0}(173,2556)(213,2556){1}
wire w30;    //: /sn:0 {0}(373,2194)(104,2194)(104,-91)(77,-91){1}
wire w123;    //: /sn:0 {0}(1269,1040)(1586,1040)(1586,974)(1654,974){1}
wire w59;    //: /sn:0 {0}(366,2527)(366,2542){1}
wire w85;    //: /sn:0 {0}(1269,880)(1540,880)(1540,894)(1654,894){1}
wire w62;    //: /sn:0 {0}(1269,790)(1616,790)(1616,849)(1654,849){1}
wire w185;    //: /sn:0 {0}(404,1170)(404,1155)(410,1155)(410,1144){1}
wire w197;    //: /sn:0 {0}(436,1343)(436,1335)(425,1335)(425,1325){1}
wire w137;    //: /sn:0 {0}(417,661)(417,650)(408,650)(408,634){1}
wire w11;    //: /sn:0 {0}(375,594)(182,594)(182,-281)(77,-281){1}
wire w57;    //: /sn:0 {0}(384,1790)(288,1790)(288,848)(-284,848){1}
wire w136;    //: /sn:0 {0}(1028,1040)(985,1040)(985,243)(458,243){1}
wire w173;    //: /sn:0 {0}(401,999)(401,986)(406,986)(406,975){1}
wire w70;    //: /sn:0 {0}(1269,830)(1584,830)(1584,869)(1654,869){1}
wire w193;    //: /sn:0 {0}(409,1839)(409,1826)(417,1826)(417,1815){1}
wire w110;    //: /sn:0 {0}(368,-361)(440,-361)(440,-391)(509,-391){1}
wire w105;    //: /sn:0 {0}(330,-312)(362,-312){1}
wire w94;    //: /sn:0 {0}(1654,919)(1524,919)(1524,930)(1269,930){1}
wire w88;    //: /sn:0 {0}(1269,900)(1523,900)(1523,904)(1654,904){1}
wire w72;    //: /sn:0 {0}(1269,840)(1577,840)(1577,874)(1654,874){1}
wire w13;    //: /sn:0 {0}(395,766)(172,766)(172,-261)(77,-261){1}
wire w5;    //: /sn:0 {0}(77,-341)(209,-341)(209,49)(367,49){1}
wire w33;    //: /sn:0 {0}(347,-376)(307,-376){1}
//: {2}(303,-376)(129,-376)(129,-326){3}
//: {4}(131,-324)(226,-324){5}
//: {6}(230,-324)(259,-324)(259,-319)(288,-319){7}
//: {8}(228,-322)(228,-301)(240,-301){9}
//: {10}(127,-324)(97,-324)(97,-426)(-260,-426)(-260,608)(-284,608){11}
//: {12}(305,-374)(305,-359)(347,-359){13}
wire w191;    //: /sn:0 {0}(424,1263)(424,1243)(405,1243)(405,1232){1}
wire w131;    //: /sn:0 {0}(1269,1080)(1639,1080)(1639,994)(1654,994){1}
wire w143;    //: /sn:0 {0}(404,481)(404,470)(393,470)(393,464)(404,464)(404,455){1}
wire w79;    //: /sn:0 {0}(1269,860)(1560,860)(1560,884)(1654,884){1}
wire w9;    //: /sn:0 {0}(77,-301)(191,-301)(191,415)(371,415){1}
wire w55;    //: /sn:0 {0}(255,2545)(317,2545)(317,2503)(332,2503){1}
wire w39;    //: /sn:0 {0}(234,2527)(234,2452)(276,2452){1}
//: {2}(280,2452)(341,2452)(341,2359)(486,2359){3}
//: {4}(490,2359)(527,2359)(527,2337){5}
//: {6}(488,2361)(488,2384){7}
//: {8}(278,2454)(278,2571)(349,2571)(349,2607){9}
wire w26;    //: /sn:0 {0}(377,1861)(118,1861)(118,-131)(77,-131){1}
//: enddecls

  //: OUT g4 (Sa) @(1322,1135) /sn:0 /w:[ 3 ]
  ALU1bit g8 (.AcarreoE(w104), .C(C), .A(w112), .B(w109), .AcarreoS(w113), .Sa(w67));   //: @(365, -256) /sz:(87, 60) /sn:0 /p:[ Ti0>1 Ti1>67 Li0>1 Li1>0 Bo0<0 Ro0<1 ]
  //: GROUND g140 (w54) @(476,-308) /sn:0 /w:[ 0 ]
  //: comment g58 @(360,1750) /sn:0
  //: /line:"24"
  //: /end
  //: comment g55 @(333,2005) /sn:0
  //: /line:"27"
  //: /end
  ALU1bit g37 (.C(C), .AcarreoE(w179), .B(w184), .A(w17), .AcarreoS(w185), .Sa(w82));   //: @(378, 1083) /sz:(87, 60) /sn:0 /p:[ Ti0>97 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<1 ]
  //: joint g13 (w0) @(325, -364) /w:[ 2 4 -1 1 ]
  //: OUT g139 (Cero) @(1738,915) /sn:0 /w:[ 0 ]
  //: joint g112 (w80) @(95, 2538) /w:[ 3 -1 4 12 ]
  //: joint g76 (C) @(716, 990) /w:[ -1 32 94 31 ]
  //: joint g111 (w32) @(295, 2481) /w:[ 1 -1 2 12 ]
  //: IN g1 (B) @(-655,763) /sn:0 /w:[ 0 ]
  //: joint g64 (C) @(717, -82) /w:[ -1 56 70 55 ]
  //: joint g11 (w0) @(325, -381) /w:[ 6 -1 8 5 ]
  //: comment g130 @(363,1155) /sn:0
  //: /line:"17"
  //: /end
  //: comment g121 @(362,385) /sn:0
  //: /line:"8"
  //: /end
  ALU1bit g50 (.C(C), .AcarreoE(w233), .B(w238), .A(w30), .AcarreoS(w239), .Sa(w240));   //: @(374, 2173) /sz:(87, 60) /sn:0 /p:[ Ti0>123 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<1 ]
  ALU1bit g28 (.C(C), .AcarreoE(w135), .B(w140), .A(w8), .AcarreoS(w141), .Sa(w73));   //: @(371, 300) /sz:(87, 60) /sn:0 /p:[ Ti0>79 Ti1>0 Li0>0 Li1>1 Bo0<0 Ro0<1 ]
  //: comment g132 @(390,1335) /sn:0
  //: /line:"19"
  //: /end
  Mux1 g19 (.C(w2), .E0(w33), .E1(w98), .Sal(w105));   //: @(289, -329) /sz:(40, 40) /sn:0 /p:[ Ti0>9 Li0>7 Li1>0 Ro0<0 ]
  //: comment g113 @(345,-295) /sn:0
  //: /line:"0"
  //: /end
  ALU1bit g38 (.C(C), .AcarreoE(w185), .B(w190), .A(w18), .AcarreoS(w191), .Sa(w192));   //: @(373, 1171) /sz:(87, 60) /sn:0 /p:[ Ti0>99 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<0 ]
  Suma g6 (.AcarreoE(w2), .B(w105), .A(w0), .AcarreoS(w104), .Suma(w100));   //: @(363, -349) /sz:(67, 60) /sn:0 /p:[ Ti0>0 Li0>1 Li1>0 Bo0<0 Ro0<0 ]
  //: comment g115 @(355,-172) /sn:0
  //: /line:"2"
  //: /end
  //: comment g53 @(339,2178) /sn:0
  //: /line:"29"
  //: /end
  Mux3 g7 (.C0(w103), .C1(w102), .C2(w2), .E0(w111), .E1(w110), .E2(w100), .E3(w54), .E4(w54), .E5(w54), .E6(w100), .E7(w65), .Sal(w66));   //: @(510, -410) /sz:(52, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>7 Li0>1 Li1>1 Li2>5 Li3>5 Li4>3 Li5>7 Li6>3 Li7>13 Ro0<0 ]
  //: joint g75 (C) @(716, 896) /w:[ -1 34 92 33 ]
  //: comment g135 @(392,2437) /sn:0
  //: /line:"31"
  //: /end
  ALU1bit g31 (.C(C), .AcarreoE(w147), .B(w133), .A(w11), .AcarreoS(w137), .Sa(w76));   //: @(376, 573) /sz:(87, 60) /sn:0 /p:[ Ti0>85 Ti1>0 Li0>1 Li1>0 Bo0<1 Ro0<1 ]
  //: joint g20 (w2) @(396, -464) /w:[ 2 -1 8 1 ]
  //: comment g124 @(375,658) /sn:0
  //: /line:"11"
  //: /end
  ALU1bit g39 (.C(C), .AcarreoE(w191), .B(w51), .A(w19), .AcarreoS(w197), .Sa(w84));   //: @(393, 1264) /sz:(87, 60) /sn:0 /p:[ Ti0>101 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<1 ]
  //: joint g68 (C) @(716, 282) /w:[ -1 48 78 47 ]
  ALU1bit g48 (.C(C), .AcarreoE(w221), .B(w226), .A(w28), .AcarreoS(w227), .Sa(w228));   //: @(363, 2006) /sz:(87, 60) /sn:0 /p:[ Ti0>119 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<1 ]
  ALU1bit g29 (.C(C), .AcarreoE(w143), .B(w42), .A(w10), .AcarreoS(w147), .Sa(w75));   //: @(373, 482) /sz:(87, 60) /sn:0 /p:[ Ti0>83 Ti1>0 Li0>1 Li1>0 Bo0<1 Ro0<1 ]
  ALU1bit g25 (.C(C), .AcarreoE(w125), .B(w37), .A(w5), .AcarreoS(w119), .Sa(w124));   //: @(368, 28) /sz:(87, 60) /sn:0 /p:[ Ti0>73 Ti1>1 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  assign {w2, w102, w103} = C; //: CONCAT g17  @(541,-514) /sn:0 /R:1 /w:[ 5 0 0 65 ] /dr:0 /tp:0 /drp:0
  //: joint g106 (w80) @(-18, 2410) /w:[ 6 8 10 5 ]
  //: comment g52 @(370,2262) /sn:0
  //: /line:"30"
  //: /end
  Overflow g107 (.A31(w32), .B31(w80), .R(w39), .SiSa(w65), .Sa(Overflow));   //: @(329, 2608) /sz:(111, 43) /sn:0 /p:[ Ti0>13 Ti1>13 Ti2>9 Ti3>11 Bo0<0 ]
  //: joint g83 (C) @(716, 1573) /w:[ -1 18 108 17 ]
  //: joint g100 (w39) @(488, 2359) /w:[ 4 -1 3 6 ]
  _GGNBUF #(2) g14 (.I(w33), .Z(w98));   //: @(246,-301) /sn:0 /w:[ 9 1 ]
  ALU1bit g47 (.C(C), .AcarreoE(w211), .B(w220), .A(w27), .AcarreoS(w221), .Sa(w92));   //: @(376, 1921) /sz:(87, 60) /sn:0 /p:[ Ti0>117 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<1 ]
  ALU1bit g44 (.C(C), .AcarreoE(w157), .B(w56), .A(w24), .AcarreoS(w175), .Sa(w89));   //: @(373, 1674) /sz:(87, 60) /sn:0 /p:[ Ti0>111 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<0 ]
  //: joint g80 (C) @(716, 1338) /w:[ -1 24 102 23 ]
  _GGAND2 #(6) g94 (.I0(w32), .I1(w80), .Z(w40));   //: @(303,2398) /sn:0 /w:[ 9 11 0 ]
  //: joint g105 (w80) @(140, 2538) /w:[ 1 -1 2 14 ]
  //: joint g21 (w33) @(129, -324) /w:[ 4 3 10 -1 ]
  //: joint g84 (C) @(716, 1659) /w:[ -1 16 110 15 ]
  //: joint g141 (w54) @(476, -363) /w:[ 2 4 6 1 ]
  ALU1bit g41 (.C(C), .AcarreoE(w203), .B(w53), .A(w21), .AcarreoS(w209), .Sa(w86));   //: @(388, 1425) /sz:(87, 60) /sn:0 /p:[ Ti0>105 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  ALU1bit g23 (.AcarreoE(w113), .C(C), .A(w3), .B(w35), .AcarreoS(w122), .Sa(w120));   //: @(366, -159) /sz:(87, 60) /sn:0 /p:[ Ti0>1 Ti1>69 Li0>1 Li1>0 Bo0<0 Ro0<1 ]
  //: comment g54 @(344,2094) /sn:0
  //: /line:"28"
  //: /end
  ALU1bit g40 (.C(C), .AcarreoE(w197), .B(w202), .A(w20), .AcarreoS(w203), .Sa(w204));   //: @(405, 1344) /sz:(87, 60) /sn:0 /p:[ Ti0>103 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  Mux1 g93 (.C(w39), .E1(w68), .E0(w80), .Sal(w55));   //: @(214, 2528) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Li0>1 Li1>0 Ro0<0 ]
  //: comment g116 @(356,-74) /sn:0
  //: /line:"3"
  //: /end
  //: comment g123 @(363,565) /sn:0
  //: /line:"10"
  //: /end
  ALU1bit g46 (.C(C), .AcarreoE(w193), .B(w207), .A(w26), .AcarreoS(w211), .Sa(w91));   //: @(378, 1840) /sz:(87, 60) /sn:0 /p:[ Ti0>115 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<0 ]
  ALU1bit g26 (.C(C), .AcarreoE(w119), .B(w38), .A(w6), .AcarreoS(w129), .Sa(w71));   //: @(369, 119) /sz:(87, 60) /sn:0 /p:[ Ti0>75 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  //: IN g0 (A) @(-135,-78) /sn:0 /w:[ 0 ]
  //: joint g90 (C) @(716, 2167) /w:[ -1 4 122 3 ]
  //: joint g82 (C) @(716, 1487) /w:[ -1 20 106 19 ]
  assign {w131, w130, w128, w127, w123, w121, w118, w117, w116, w115, w114, w101, w99, w97, w95, w94, w93, w90, w88, w87, w85, w83, w79, w77, w72, w70, w69, w64, w63, w62, w50, w43} = Sa; //: CONCAT g136  @(1264,925) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /dr:0 /tp:0 /drp:0
  //: comment g128 @(364,983) /sn:0
  //: /line:"15"
  //: /end
  ALU1bit g33 (.C(C), .AcarreoE(w155), .B(w45), .A(w13), .AcarreoS(w161), .Sa(w78));   //: @(396, 745) /sz:(87, 60) /sn:0 /p:[ Ti0>89 Ti1>0 Li0>1 Li1>0 Bo0<1 Ro0<1 ]
  Mux3 g91 (.C2(w39), .C1(w34), .C0(w1), .E7(w49), .E6(w65), .E5(w49), .E4(w49), .E3(w49), .E2(w65), .E1(w41), .E0(w40), .Sal(w52));   //: @(468, 2385) /sz:(52, 85) /sn:0 /p:[ Ti0>7 Ti1>1 Ti2>1 Li0>11 Li1>0 Li2>7 Li3>0 Li4>3 Li5>5 Li6>1 Li7>1 Ro0<1 ]
  ALU1bit g49 (.C(C), .AcarreoE(w227), .B(w61), .A(w29), .AcarreoS(w233), .Sa(w234));   //: @(388, 2094) /sz:(87, 60) /sn:0 /p:[ Ti0>121 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<1 ]
  _GGNOR32 #(64) g137 (.I0(w43), .I1(w50), .I2(w62), .I3(w63), .I4(w64), .I5(w69), .I6(w70), .I7(w72), .I8(w77), .I9(w79), .I10(w83), .I11(w85), .I12(w87), .I13(w88), .I14(w90), .I15(w93), .I16(w94), .I17(w95), .I18(w97), .I19(w99), .I20(w101), .I21(w114), .I22(w115), .I23(w116), .I24(w117), .I25(w118), .I26(w121), .I27(w123), .I28(w127), .I29(w128), .I30(w130), .I31(w131), .Z(Cero));   //: @(1665,916) /sn:0 /w:[ 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ]
  //: joint g61 (C) @(573, -536) /w:[ 61 62 -1 64 ]
  ALU1bit g51 (.C(C), .AcarreoE(w239), .B(w244), .A(w31), .AcarreoS(w245), .Sa(w96));   //: @(395, 2257) /sz:(87, 60) /sn:0 /p:[ Ti0>125 Ti1>0 Li0>0 Li1>0 Bo0<0 Ro0<1 ]
  ALU1bit g34 (.C(C), .AcarreoE(w161), .B(w166), .A(w14), .AcarreoS(w167), .Sa(w168));   //: @(378, 830) /sz:(87, 60) /sn:0 /p:[ Ti0>91 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  assign {w80, w244, w238, w61, w226, w220, w207, w57, w56, w151, w214, w53, w202, w51, w190, w184, w178, w172, w166, w45, w44, w133, w42, w152, w140, w134, w38, w37, w36, w35, w109, w33} = B; //: CONCAT g3  @(-289,763) /sn:0 /R:2 /w:[ 9 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1 11 1 ] /dr:0 /tp:0 /drp:0
  //: joint g86 (C) @(716, 1826) /w:[ -1 12 114 11 ]
  //: joint g89 (C) @(716, 2077) /w:[ -1 6 120 5 ]
  assign {w32, w31, w30, w29, w28, w27, w26, w25, w24, w23, w22, w21, w20, w19, w18, w17, w16, w15, w14, w13, w12, w11, w10, w9, w8, w7, w6, w5, w4, w3, w112, w0} = A; //: CONCAT g2  @(72,-226) /sn:0 /R:2 /w:[ 11 1 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 9 1 ] /dr:0 /tp:0 /drp:0
  //: joint g65 (C) @(717, 4) /w:[ -1 54 72 53 ]
  //: joint g77 (C) @(716, 1092) /w:[ -1 30 96 29 ]
  //: joint g110 (w65) @(424, 2494) /w:[ -1 7 8 10 ]
  //: comment g59 @(355,1673) /sn:0
  //: /line:"23"
  //: /end
  //: joint g72 (C) @(716, 655) /w:[ -1 40 86 39 ]
  assign {w39, w34, w1} = C; //: CONCAT g98  @(537,2332) /sn:0 /R:1 /w:[ 5 0 0 0 ] /dr:0 /tp:0 /drp:0
  //: joint g99 (C) @(537, 2251) /w:[ 2 -1 124 1 ]
  //: IN g16 (C) @(541,-548) /sn:0 /R:3 /w:[ 63 ]
  //: joint g96 (w65) @(424, 2453) /w:[ 3 4 -1 6 ]
  //: joint g103 (w32) @(98, 2392) /w:[ 8 10 -1 7 ]
  //: comment g122 @(363,473) /sn:0
  //: /line:"9"
  //: /end
  _GGOR2 #(6) g10 (.I0(w0), .I1(w33), .Z(w110));   //: @(358,-361) /sn:0 /w:[ 3 13 0 ]
  //: joint g78 (C) @(716, 1149) /w:[ -1 28 98 27 ]
  //: joint g87 (C) @(716, 1911) /w:[ -1 10 116 9 ]
  //: comment g129 @(364,1074) /sn:0
  //: /line:"16"
  //: /end
  ALU1bit g32 (.C(C), .AcarreoE(w137), .B(w44), .A(w12), .AcarreoS(w155), .Sa(w156));   //: @(386, 662) /sz:(87, 60) /sn:0 /p:[ Ti0>87 Ti1>0 Li0>1 Li1>0 Bo0<1 Ro0<1 ]
  ALU1bit g27 (.C(C), .AcarreoE(w129), .B(w134), .A(w7), .AcarreoS(w135), .Sa(w136));   //: @(370, 212) /sz:(87, 60) /sn:0 /p:[ Ti0>77 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  //: joint g102 (w65) @(446, 2453) /w:[ 1 -1 2 12 ]
  //: joint g143 (w49) @(451, 2446) /w:[ -1 6 5 8 ]
  //: joint g69 (C) @(716, 371) /w:[ -1 46 80 45 ]
  //: comment g57 @(344,1839) /sn:0
  //: /line:"25"
  //: /end
  _GGAND2 #(6) g9 (.I0(w0), .I1(w33), .Z(w111));   //: @(358,-378) /sn:0 /w:[ 7 0 0 ]
  //: comment g119 @(357,206) /sn:0
  //: /line:"6"
  //: /end
  //: joint g142 (w49) @(451, 2463) /w:[ 10 9 -1 12 ]
  //: joint g15 (w100) @(455, -342) /w:[ 2 4 -1 1 ]
  //: joint g71 (C) @(716, 559) /w:[ -1 42 84 41 ]
  //: comment g131 @(379,1252) /sn:0
  //: /line:"18"
  //: /end
  //: joint g67 (C) @(716, 195) /w:[ -1 50 76 49 ]
  //: comment g127 @(365,901) /sn:0
  //: /line:"14"
  //: /end
  ALU1bit g43 (.C(C), .AcarreoE(w215), .B(w151), .A(w23), .AcarreoS(w157), .Sa(w159));   //: @(378, 1593) /sz:(87, 60) /sn:0 /p:[ Ti0>109 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<0 ]
  //: joint g104 (w32) @(98, 2407) /w:[ 4 6 -1 3 ]
  //: joint g62 (C) @(717, -279) /w:[ -1 60 66 59 ]
  //: joint g73 (C) @(716, 739) /w:[ -1 38 88 37 ]
  //: joint g88 (C) @(716, 1996) /w:[ -1 8 118 7 ]
  //: joint g138 (Sa) @(1138, 1135) /w:[ 2 1 4 -1 ]
  ALU1bit g42 (.C(C), .AcarreoE(w209), .B(w214), .A(w22), .AcarreoS(w215), .Sa(w216));   //: @(385, 1508) /sz:(87, 60) /sn:0 /p:[ Ti0>107 Ti1>0 Li0>0 Li1>0 Bo0<1 Ro0<0 ]
  //: joint g63 (C) @(717, -174) /w:[ -1 58 68 57 ]
  //: joint g74 (C) @(716, 824) /w:[ -1 36 90 35 ]
  //: joint g109 (w39) @(278, 2452) /w:[ 2 -1 1 8 ]
  //: comment g133 @(374,1410) /sn:0
  //: /line:"20"
  //: /end
  //: comment g56 @(346,1923) /sn:0
  //: /line:"26"
  //: /end
  assign Sa = {w52, w96, w240, w234, w228, w92, w91, w195, w89, w159, w216, w86, w204, w84, w192, w82, w81, w174, w168, w78, w156, w76, w75, w74, w73, w136, w71, w124, w126, w120, w67, w66}; //: CONCAT g5  @(1033,1135) /sn:0 /w:[ 5 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:1 /tp:0 /drp:1
  //: joint g79 (C) @(716, 1236) /w:[ -1 26 100 25 ]
  _GGOR2 #(6) g95 (.I0(w32), .I1(w80), .Z(w41));   //: @(303,2415) /sn:0 /w:[ 5 7 0 ]
  //: comment g117 @(350,27) /sn:0
  //: /line:"4"
  //: /end
  ALU1bit g36 (.C(C), .AcarreoE(w173), .B(w178), .A(w16), .AcarreoS(w179), .Sa(w81));   //: @(370, 1000) /sz:(87, 60) /sn:0 /p:[ Ti0>95 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  ALU1bit g24 (.AcarreoE(w122), .C(C), .A(w4), .B(w36), .AcarreoS(w125), .Sa(w126));   //: @(367, -62) /sz:(87, 60) /sn:0 /p:[ Ti0>1 Ti1>71 Li0>1 Li1>0 Bo0<0 Ro0<1 ]
  //: joint g85 (C) @(716, 1746) /w:[ -1 14 112 13 ]
  Suma g92 (.AcarreoE(w245), .A(w32), .B(w55), .AcarreoS(w59), .Suma(w65));   //: @(333, 2466) /sz:(67, 60) /sn:0 /p:[ Ti0>1 Li0>0 Li1>1 Bo0<0 Ro0<9 ]
  //: joint g144 (w49) @(439, 2432) /w:[ 1 2 -1 4 ]
  //: comment g125 @(380,735) /sn:0
  //: /line:"12"
  //: /end
  //: comment g60 @(360,1587) /sn:0
  //: /line:"22"
  //: /end
  //: joint g81 (C) @(716, 1414) /w:[ -1 22 104 21 ]
  _GGNBUF #(2) g101 (.I(w80), .Z(w68));   //: @(163,2556) /sn:0 /w:[ 15 0 ]
  ALU1bit g35 (.C(C), .AcarreoE(w167), .B(w172), .A(w15), .AcarreoS(w173), .Sa(w174));   //: @(374, 914) /sz:(87, 60) /sn:0 /p:[ Ti0>93 Ti1>0 Li0>1 Li1>0 Bo0<1 Ro0<1 ]
  //: joint g22 (w33) @(228, -324) /w:[ 6 -1 5 8 ]
  //: joint g70 (C) @(716, 459) /w:[ -1 44 82 43 ]
  //: comment g126 @(375,809) /sn:0
  //: /line:"13"
  //: /end
  ALU1bit g45 (.C(C), .AcarreoE(w175), .B(w57), .A(w25), .AcarreoS(w193), .Sa(w195));   //: @(385, 1754) /sz:(87, 60) /sn:0 /p:[ Ti0>113 Ti1>0 Li0>0 Li1>1 Bo0<1 Ro0<0 ]
  //: joint g66 (C) @(717, 104) /w:[ -1 52 74 51 ]
  //: GROUND g97 (w49) @(451,2504) /sn:0 /w:[ 13 ]
  //: comment g114 @(353,-261) /sn:0
  //: /line:"1"
  //: /end
  //: comment g120 @(356,294) /sn:0
  //: /line:"7"
  //: /end
  //: joint g18 (w2) @(530, -464) /w:[ -1 4 3 6 ]
  //: joint g12 (w33) @(305, -376) /w:[ 1 -1 2 12 ]
  ALU1bit g30 (.C(C), .AcarreoE(w141), .B(w152), .A(w9), .AcarreoS(w143), .Sa(w74));   //: @(372, 394) /sz:(87, 60) /sn:0 /p:[ Ti0>81 Ti1>1 Li0>0 Li1>1 Bo0<1 Ro0<1 ]
  //: OUT g108 (Overflow) @(410,2708) /sn:0 /w:[ 1 ]
  //: comment g134 @(371,1496) /sn:0
  //: /line:"21"
  //: /end
  //: comment g118 @(351,115) /sn:0
  //: /line:"5"
  //: /end

endmodule
//: /netlistEnd

//: /netlistBegin Mux3
module Mux3(E0, E4, C0, C1, C2, E7, E6, E2, E3, E5, E1, Sal);
//: interface  /sz:(52, 85) /bd:[ Ti0>C0(42/52) Ti1>C1(31/52) Ti2>C2(20/52) Li0>E0(7/85) Li1>E1(19/85) Li2>E2(27/85) Li3>E3(38/85) Li4>E4(47/85) Li5>E5(57/85) Li6>E6(68/85) Li7>E7(78/85) Ro0<Sal(41/85) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input E7;    //: /sn:0 {0}(502,399)(292,399)(292,410)(277,410){1}
input C0;    //: /sn:0 {0}(422,116)(422,174){1}
//: {2}(424,176)(501,176){3}
//: {4}(422,178)(422,202){5}
//: {6}(424,204)(502,204){7}
//: {8}(422,206)(422,232){9}
//: {10}(424,234)(502,234){11}
//: {12}(422,236)(422,264){13}
//: {14}(424,266)(434,266)(434,267)(502,267){15}
//: {16}(422,268)(422,300){17}
//: {18}(424,302)(434,302)(434,301)(503,301){19}
//: {20}(422,304)(422,333){21}
//: {22}(424,335)(434,335)(434,336)(503,336){23}
//: {24}(422,337)(422,367){25}
//: {26}(424,369)(434,369)(434,370)(503,370){27}
//: {28}(422,371)(422,404)(502,404){29}
input E1;    //: /sn:0 {0}(502,199)(288,199)(288,213)(273,213){1}
input E2;    //: /sn:0 {0}(502,229)(290,229)(290,248)(275,248){1}
input E0;    //: /sn:0 {0}(501,171)(287,171)(287,180)(272,180){1}
input C2;    //: /sn:0 {0}(501,186)(389,186)(389,184)(379,184){1}
//: {2}(377,182)(377,116){3}
//: {4}(377,186)(377,211){5}
//: {6}(379,213)(389,213)(389,214)(502,214){7}
//: {8}(377,215)(377,243){9}
//: {10}(379,245)(389,245)(389,244)(502,244){11}
//: {12}(377,247)(377,275){13}
//: {14}(379,277)(502,277){15}
//: {16}(377,279)(377,310){17}
//: {18}(379,312)(389,312)(389,311)(503,311){19}
//: {20}(377,314)(377,342){21}
//: {22}(379,344)(389,344)(389,346)(503,346){23}
//: {24}(377,346)(377,376){25}
//: {26}(379,378)(389,378)(389,380)(503,380){27}
//: {28}(377,380)(377,412)(389,412)(389,414)(502,414){29}
output Sal;    //: /sn:0 {0}(639,287)(731,287)(731,291)(741,291){1}
input E4;    //: /sn:0 {0}(503,296)(286,296)(286,314)(271,314){1}
input E3;    //: /sn:0 {0}(502,262)(288,262)(288,277)(273,277){1}
input E5;    //: /sn:0 {0}(503,331)(288,331)(288,349)(273,349){1}
input C1;    //: /sn:0 {0}(503,375)(410,375)(410,373)(400,373){1}
//: {2}(398,371)(398,344){3}
//: {4}(400,342)(410,342)(410,341)(503,341){5}
//: {6}(398,340)(398,305){7}
//: {8}(400,303)(410,303)(410,306)(503,306){9}
//: {10}(398,301)(398,272){11}
//: {12}(400,270)(410,270)(410,272)(502,272){13}
//: {14}(398,268)(398,238){15}
//: {16}(400,236)(410,236)(410,239)(502,239){17}
//: {18}(398,234)(398,211){19}
//: {20}(400,209)(502,209){21}
//: {22}(398,207)(398,181){23}
//: {24}(400,179)(410,179)(410,181)(501,181){25}
//: {26}(398,177)(398,116){27}
//: {28}(398,375)(398,409)(502,409){29}
input E6;    //: /sn:0 {0}(503,365)(291,365)(291,378)(276,378){1}
wire w14;    //: /sn:0 {0}(524,303)(583,303)(583,290)(618,290){1}
wire w20;    //: /sn:0 {0}(524,372)(597,372)(597,300)(618,300){1}
wire w23;    //: /sn:0 {0}(523,406)(603,406)(603,305)(618,305){1}
wire w8;    //: /sn:0 {0}(523,236)(589,236)(589,280)(618,280){1}
wire w17;    //: /sn:0 {0}(524,338)(591,338)(591,295)(618,295){1}
wire w2;    //: /sn:0 {0}(522,178)(603,178)(603,270)(618,270){1}
wire w11;    //: /sn:0 {0}(523,269)(584,269)(584,285)(618,285){1}
wire w5;    //: /sn:0 {0}(523,206)(596,206)(596,275)(618,275){1}
//: enddecls

  //: IN g4 (E0) @(270,180) /sn:0 /w:[ 1 ]
  //: IN g8 (E4) @(269,314) /sn:0 /w:[ 1 ]
  //: IN g3 (C0) @(422,114) /sn:0 /R:3 /w:[ 0 ]
  _GGAND4 #(10) g13 (.I0(E1), .I1(C0), .I2(!C1), .I3(!C2), .Z(w5));   //: @(513,206) /sn:0 /w:[ 0 7 21 7 0 ]
  //: joint g34 (C1) @(398, 342) /w:[ 4 6 -1 3 ]
  //: IN g2 (C1) @(398,114) /sn:0 /R:3 /w:[ 27 ]
  //: IN g1 (C2) @(377,114) /sn:0 /R:3 /w:[ 3 ]
  //: IN g11 (E7) @(275,410) /sn:0 /w:[ 1 ]
  _GGAND4 #(10) g16 (.I0(E4), .I1(!C0), .I2(!C1), .I3(C2), .Z(w14));   //: @(514,303) /sn:0 /w:[ 0 19 9 19 0 ]
  //: IN g10 (E6) @(274,378) /sn:0 /w:[ 1 ]
  _GGAND4 #(10) g19 (.I0(E7), .I1(C0), .I2(C1), .I3(C2), .Z(w23));   //: @(513,406) /sn:0 /w:[ 0 29 29 29 0 ]
  //: joint g27 (C0) @(422, 369) /w:[ 26 25 -1 28 ]
  //: joint g32 (C1) @(398, 270) /w:[ 12 14 -1 11 ]
  //: IN g6 (E2) @(273,248) /sn:0 /w:[ 1 ]
  //: joint g38 (C2) @(377, 378) /w:[ 26 25 -1 28 ]
  //: IN g7 (E3) @(271,277) /sn:0 /w:[ 1 ]
  //: IN g9 (E5) @(271,349) /sn:0 /w:[ 1 ]
  _GGAND4 #(10) g15 (.I0(E3), .I1(C0), .I2(C1), .I3(!C2), .Z(w11));   //: @(513,269) /sn:0 /w:[ 0 15 13 15 0 ]
  _GGOR8 #(18) g20 (.I0(w2), .I1(w5), .I2(w8), .I3(w11), .I4(w14), .I5(w17), .I6(w20), .I7(w23), .Z(Sal));   //: @(629,287) /sn:0 /w:[ 1 1 1 1 1 1 1 1 0 ]
  //: joint g31 (C1) @(398, 236) /w:[ 16 18 -1 15 ]
  //: joint g39 (C2) @(377, 344) /w:[ 22 21 -1 24 ]
  //: joint g43 (C2) @(377, 213) /w:[ 6 5 -1 8 ]
  _GGAND4 #(10) g17 (.I0(E5), .I1(C0), .I2(!C1), .I3(C2), .Z(w17));   //: @(514,338) /sn:0 /w:[ 0 23 5 23 0 ]
  //: joint g25 (C0) @(422, 302) /w:[ 18 17 -1 20 ]
  //: joint g29 (C1) @(398, 179) /w:[ 24 26 -1 23 ]
  //: joint g42 (C2) @(377, 245) /w:[ 10 9 -1 12 ]
  //: IN g5 (E1) @(271,213) /sn:0 /w:[ 1 ]
  _GGAND4 #(10) g14 (.I0(E2), .I1(!C0), .I2(C1), .I3(!C2), .Z(w8));   //: @(513,236) /sn:0 /w:[ 0 11 17 11 0 ]
  //: joint g44 (C2) @(377, 184) /w:[ 1 2 -1 4 ]
  //: joint g21 (C0) @(422, 176) /w:[ 2 1 -1 4 ]
  //: joint g24 (C0) @(422, 266) /w:[ 14 13 -1 16 ]
  //: joint g23 (C0) @(422, 234) /w:[ 10 9 -1 12 ]
  //: joint g41 (C2) @(377, 277) /w:[ 14 13 -1 16 ]
  //: joint g40 (C2) @(377, 312) /w:[ 18 17 -1 20 ]
  //: OUT g0 (Sal) @(738,291) /sn:0 /w:[ 1 ]
  //: joint g22 (C0) @(422, 204) /w:[ 6 5 -1 8 ]
  //: joint g26 (C0) @(422, 335) /w:[ 22 21 -1 24 ]
  //: joint g35 (C1) @(398, 373) /w:[ 1 2 -1 28 ]
  _GGAND4 #(10) g12 (.I0(E0), .I1(!C0), .I2(!C1), .I3(!C2), .Z(w2));   //: @(512,178) /sn:0 /w:[ 0 3 25 0 0 ]
  _GGAND4 #(10) g18 (.I0(E6), .I1(!C0), .I2(C1), .I3(C2), .Z(w20));   //: @(514,372) /sn:0 /w:[ 0 27 0 27 0 ]
  //: joint g30 (C1) @(398, 209) /w:[ 20 22 -1 19 ]
  //: joint g33 (C1) @(398, 303) /w:[ 8 10 -1 7 ]

endmodule
//: /netlistEnd

//: /netlistBegin Overflow
module Overflow(Sa, SiSa, B31, A31, R);
//: interface  /sz:(111, 43) /bd:[ Ti0>SiSa(85/111) Ti1>R(20/111) Ti2>B31(63/111) Ti3>A31(42/111) Bo0<Sa(54/111) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input A31;    //: /sn:0 {0}(286,245)(286,113){1}
//: {2}(288,111)(334,111){3}
//: {4}(338,111)(383,111){5}
//: {6}(387,111)(427,111)(427,244){7}
//: {8}(385,113)(385,245){9}
//: {10}(336,113)(336,123)(337,123)(337,246){11}
//: {12}(284,111)(130,111){13}
input SiSa;    //: /sn:0 {0}(126,190)(294,190){1}
//: {2}(298,190)(345,190){3}
//: {4}(349,190)(393,190){5}
//: {6}(397,190)(437,190)(437,244){7}
//: {8}(395,192)(395,245){9}
//: {10}(347,192)(347,246){11}
//: {12}(296,192)(296,245){13}
input R;    //: /sn:0 {0}(281,245)(281,88)(280,88)(280,78){1}
//: {2}(282,76)(327,76){3}
//: {4}(331,76)(378,76){5}
//: {6}(382,76)(422,76)(422,244){7}
//: {8}(380,78)(380,245){9}
//: {10}(329,78)(329,88)(332,88)(332,246){11}
//: {12}(278,76)(127,76){13}
output Sa;    //: /sn:0 {0}(616,416)(364,416)(364,353){1}
input B31;    //: /sn:0 {0}(126,152)(251,152)(251,151)(290,151){1}
//: {2}(294,151)(339,151){3}
//: {4}(343,151)(387,151){5}
//: {6}(391,151)(432,151)(432,244){7}
//: {8}(389,153)(389,163)(390,163)(390,245){9}
//: {10}(341,153)(341,163)(342,163)(342,246){11}
//: {12}(292,153)(292,163)(291,163)(291,245){13}
wire w2;    //: /sn:0 {0}(361,332)(361,277)(340,277)(340,267){1}
wire w12;    //: /sn:0 {0}(289,266)(289,317)(356,317)(356,332){1}
wire w11;    //: /sn:0 {0}(430,265)(430,317)(371,317)(371,332){1}
wire w5;    //: /sn:0 {0}(366,332)(366,276)(388,276)(388,266){1}
//: enddecls

  _GGAND4 #(10) g8 (.I0(!SiSa), .I1(!B31), .I2(A31), .I3(R), .Z(w11));   //: @(430,255) /sn:0 /R:3 /w:[ 7 7 7 7 0 ]
  //: OUT g4 (Sa) @(613,416) /sn:0 /w:[ 0 ]
  //: joint g13 (R) @(380, 76) /w:[ 6 -1 5 8 ]
  //: IN g3 (SiSa) @(124,190) /sn:0 /w:[ 0 ]
  //: IN g2 (B31) @(124,152) /sn:0 /w:[ 0 ]
  //: IN g1 (A31) @(128,111) /sn:0 /w:[ 13 ]
  //: joint g16 (A31) @(336, 111) /w:[ 4 -1 3 10 ]
  //: joint g11 (B31) @(389, 151) /w:[ 6 -1 5 8 ]
  //: joint g10 (SiSa) @(395, 190) /w:[ 6 -1 5 8 ]
  //: joint g19 (B31) @(292, 151) /w:[ 2 -1 1 12 ]
  _GGAND4 #(10) g6 (.I0(!SiSa), .I1(B31), .I2(A31), .I3(!R), .Z(w2));   //: @(340,257) /sn:0 /R:3 /w:[ 11 11 11 11 1 ]
  _GGOR4 #(10) g9 (.I0(w11), .I1(w5), .I2(w2), .I3(w12), .Z(Sa));   //: @(364,343) /sn:0 /R:3 /w:[ 1 0 0 1 1 ]
  _GGAND4 #(10) g7 (.I0(SiSa), .I1(B31), .I2(!A31), .I3(R), .Z(w5));   //: @(388,256) /sn:0 /R:3 /w:[ 9 9 9 9 1 ]
  //: joint g20 (A31) @(286, 111) /w:[ 2 -1 12 1 ]
  //: joint g15 (B31) @(341, 151) /w:[ 4 -1 3 10 ]
  //: joint g17 (R) @(329, 76) /w:[ 4 -1 3 10 ]
  //: joint g14 (SiSa) @(347, 190) /w:[ 4 -1 3 10 ]
  _GGAND4 #(10) g5 (.I0(SiSa), .I1(!B31), .I2(!A31), .I3(!R), .Z(w12));   //: @(289,256) /sn:0 /R:3 /w:[ 13 13 0 0 0 ]
  //: joint g21 (R) @(280, 76) /w:[ 2 -1 12 1 ]
  //: IN g0 (R) @(125,76) /sn:0 /w:[ 13 ]
  //: joint g18 (SiSa) @(296, 190) /w:[ 2 -1 1 12 ]
  //: joint g12 (A31) @(385, 111) /w:[ 6 -1 5 8 ]

endmodule
//: /netlistEnd

//: /netlistBegin LatchD
module LatchD(Q, D, C, nQ);
//: interface  /sz:(75, 48) /bd:[ Li0>C(29/48) Li1>D(14/48) Ro0<nQ(31/48) Ro1<Q(12/48) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output Q;    //: /sn:0 {0}(339,117)(379,117){1}
//: {2}(383,117)(425,117)(425,103)(438,103){3}
//: {4}(381,119)(381,161)(313,161)(313,176)(323,176){5}
output nQ;    //: /sn:0 {0}(344,179)(388,179){1}
//: {2}(392,179)(416,179)(416,162)(429,162){3}
//: {4}(390,177)(390,132)(300,132)(300,119)(318,119){5}
input D;    //: /sn:0 {0}(86,90)(118,90){1}
//: {2}(122,90)(167,90)(167,102)(180,102){3}
//: {4}(120,92)(120,155)(181,155){5}
input C;    //: /sn:0 {0}(25,183)(106,183)(106,160)(138,160){1}
//: {2}(142,160)(181,160){3}
//: {4}(140,158)(140,107)(180,107){5}
wire w2;    //: /sn:0 {0}(201,105)(303,105)(303,114)(318,114){1}
wire w5;    //: /sn:0 {0}(202,158)(216,158)(216,194)(223,194)(223,181)(323,181){1}
//: enddecls

  //: OUT g4 (Q) @(435,103) /sn:0 /w:[ 3 ]
  //: joint g8 (D) @(120, 90) /w:[ 2 -1 1 4 ]
  _GGNOR2 #(4) g3 (.I0(Q), .I1(w5), .Z(nQ));   //: @(334,179) /sn:0 /w:[ 5 1 0 ]
  _GGNOR2 #(4) g2 (.I0(w2), .I1(nQ), .Z(Q));   //: @(329,117) /sn:0 /w:[ 1 5 0 ]
  _GGAND2 #(6) g1 (.I0(D), .I1(C), .Z(w5));   //: @(192,158) /sn:0 /w:[ 5 3 0 ]
  //: joint g11 (nQ) @(390, 179) /w:[ 2 4 1 -1 ]
  //: joint g10 (Q) @(381, 117) /w:[ 2 -1 1 4 ]
  //: IN g6 (D) @(84,90) /sn:0 /w:[ 0 ]
  //: IN g7 (C) @(23,183) /sn:0 /w:[ 0 ]
  //: joint g9 (C) @(140, 160) /w:[ 2 4 1 -1 ]
  //: OUT g5 (nQ) @(426,162) /sn:0 /w:[ 3 ]
  _GGAND2 #(6) g0 (.I0(!D), .I1(C), .Z(w2));   //: @(191,105) /sn:0 /w:[ 3 5 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin Mux1
module Mux1(Sal, E1, E0, C);
//: interface  /sz:(40, 40) /bd:[ Ti0>C(20/40) Li0>E0(10/40) Li1>E1(28/40) Ro0<Sal(17/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input E1;    //: /sn:0 {0}(293,241)(401,241){1}
input E0;    //: /sn:0 {0}(293,202)(398,202){1}
output Sal;    //: /sn:0 {0}(493,222)(537,222){1}
input C;    //: /sn:0 {0}(359,143)(359,205){1}
//: {2}(361,207)(398,207){3}
//: {4}(359,209)(359,246)(401,246){5}
wire w2;    //: /sn:0 {0}(419,205)(459,205)(459,219)(472,219){1}
wire w5;    //: /sn:0 {0}(422,244)(458,244)(458,224)(472,224){1}
//: enddecls

  _GGAND2 #(6) g4 (.I0(E0), .I1(!C), .Z(w2));   //: @(409,205) /sn:0 /w:[ 1 3 0 ]
  //: OUT g3 (Sal) @(534,222) /sn:0 /w:[ 1 ]
  //: IN g2 (E1) @(291,241) /sn:0 /w:[ 0 ]
  //: IN g1 (E0) @(291,202) /sn:0 /w:[ 0 ]
  _GGOR2 #(6) g6 (.I0(w2), .I1(w5), .Z(Sal));   //: @(483,222) /sn:0 /w:[ 1 1 0 ]
  //: joint g7 (C) @(359, 207) /w:[ 2 1 -1 4 ]
  _GGAND2 #(6) g5 (.I0(E1), .I1(C), .Z(w5));   //: @(412,244) /sn:0 /w:[ 1 5 0 ]
  //: IN g0 (C) @(359,141) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FlipFlopJK
module FlipFlopJK(Q, nQ, J, Reloj, R, K);
//: interface  /sz:(77, 58) /bd:[ Ti0>R(36/77) Li0>K(39/58) Li1>J(13/58) Bi0>Reloj(37/77) Ro0<nQ(39/58) Ro1<Q(13/58) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output nQ;    //: /sn:0 {0}(504,311)(538,311)(538,326)(549,326)(549,342)(581,342){1}
output Q;    //: /sn:0 {0}(504,284)(531,284){1}
//: {2}(535,284)(551,284)(551,268)(581,268){3}
//: {4}(533,282)(533,173)(184,173)(184,210){5}
//: {6}(186,212)(207,212){7}
//: {8}(184,214)(184,259)(207,259){9}
input K;    //: /sn:0 {0}(39,256)(95,256){1}
input R;    //: /sn:0 {0}(70,149)(70,202){1}
//: {2}(72,204)(95,204){3}
//: {4}(70,206)(70,251)(95,251){5}
input J;    //: /sn:0 {0}(95,209)(35,209){1}
supply0 w8;    //: /sn:0 {0}(645,307)(645,241){1}
//: {2}(645,237)(645,220)(653,220){3}
//: {4}(657,220)(673,220){5}
//: {6}(675,218)(675,134)(701,134){7}
//: {8}(675,222)(675,251)(690,251){9}
//: {10}(655,222)(655,256)(690,256){11}
//: {12}(643,239)(631,239)(631,129)(701,129){13}
supply1 w12;    //: /sn:0 {0}(513,367)(513,382)(445,382)(445,336){1}
input Reloj;    //: /sn:0 {0}(228,370)(364,370)(364,308)(373,308){1}
wire w6;    //: /sn:0 {0}(711,256)(813,256)(813,241)(828,241){1}
wire w7;    //: /sn:0 {0}(294,232)(358,232)(358,282)(373,282){1}
wire w14;    //: /sn:0 {0}(228,257)(258,257)(258,234)(273,234){1}
wire w4;    //: /sn:0 {0}(690,261)(680,261)(680,291)(903,291)(903,239)(892,239)(892,238)(886,238){1}
//: {2}(884,236)(884,170)(819,170)(819,156)(831,156){3}
//: {4}(882,238)(864,238)(864,239)(849,239){5}
wire w3;    //: /sn:0 {0}(852,154)(883,154)(883,155)(909,155){1}
//: {2}(911,153)(911,100)(697,100)(697,124)(701,124){3}
//: {4}(911,157)(911,222)(824,222)(824,236)(828,236){5}
wire w2;    //: /sn:0 {0}(722,129)(816,129)(816,151)(831,151){1}
wire w10;    //: /sn:0 {0}(228,210)(258,210)(258,229)(273,229){1}
wire w13;    //: /sn:0 {0}(116,254)(207,254){1}
wire w5;    //: /sn:0 {0}(116,207)(207,207){1}
//: enddecls

  //: OUT g4 (Q) @(578,268) /sn:0 /w:[ 3 ]
  _GGNOR2 #(4) g8 (.I0(w3), .I1(w6), .Z(w4));   //: @(839,239) /sn:0 /w:[ 5 1 5 ]
  //: comment g37 @(89,170) /sn:0
  //: /line:"Reset"
  //: /end
  _GGOR2 #(6) g34 (.I0(R), .I1(K), .Z(w13));   //: @(106,254) /sn:0 /w:[ 5 1 0 ]
  //: OUT g3 (nQ) @(578,342) /sn:0 /w:[ 1 ]
  //: comment g13 @(640,194) /sn:0
  //: /line:"Reloj"
  //: /end
  //: IN g2 (J) @(33,209) /sn:0 /w:[ 1 ]
  //: IN g1 (Reloj) @(226,370) /sn:0 /w:[ 0 ]
  //: joint g11 (w4) @(884, 238) /w:[ 1 2 4 -1 ]
  //: comment g16 @(906,244) /sn:0
  //: /line:"nQ"
  //: /end
  //: joint g28 (w8) @(675, 220) /w:[ -1 6 5 8 ]
  //: joint g10 (w3) @(911, 155) /w:[ -1 2 1 4 ]
  //: IN g32 (R) @(70,147) /sn:0 /R:3 /w:[ 0 ]
  //: GROUND g27 (w8) @(645,313) /sn:0 /w:[ 0 ]
  //: VDD g19 (w12) @(524,367) /sn:0 /w:[ 0 ]
  _GGAND3 #(8) g6 (.I0(w8), .I1(w8), .I2(w4), .Z(w6));   //: @(701,256) /sn:0 /w:[ 9 11 0 0 ]
  _GGNOR2 #(4) g7 (.I0(w2), .I1(w4), .Z(w3));   //: @(842,154) /sn:0 /w:[ 1 3 0 ]
  //: frame g9 @(625,45) /sn:0 /wi:337 /ht:293 /tx:""
  //: comment g31 @(374,67) /sn:0
  //: /line:"Flanco ascendente"
  //: /line:""
  //: /line:"Para iniciar poner k a 1 y J a 0"
  //: /line:"Se inicia a 0"
  //: /line:""
  //: /line:"Con poner 1 en R basta"
  //: /end
  _GGAND2 #(6) g20 (.I0(w5), .I1(!Q), .Z(w10));   //: @(218,210) /sn:0 /w:[ 1 7 0 ]
  //: comment g15 @(661,256) /sn:0
  //: /line:"J"
  //: /end
  //: joint g29 (w8) @(655, 220) /w:[ 4 -1 3 10 ]
  //: frame g25 @(156,145) /sn:0 /wi:159 /ht:135 /tx:""
  //: comment g17 @(917,149) /sn:0
  //: /line:"Q"
  //: /end
  _GGAND3 #(8) g5 (.I0(w3), .I1(w8), .I2(w8), .Z(w2));   //: @(712,129) /sn:0 /w:[ 3 13 7 0 ]
  //: comment g14 @(678,114) /sn:0
  //: /line:"K"
  //: /end
  //: frame g36 @(55,168) /sn:0 /wi:93 /ht:101 /tx:""
  //: joint g24 (Q) @(184, 212) /w:[ 6 5 -1 8 ]
  _GGAND2 #(6) g21 (.I0(!w13), .I1(Q), .Z(w14));   //: @(218,257) /sn:0 /w:[ 1 9 0 ]
  //: joint g23 (Q) @(533, 284) /w:[ 2 4 1 -1 ]
  //: joint g35 (R) @(70, 204) /w:[ 2 1 -1 4 ]
  //: comment g26 @(201,148) /sn:0
  //: /line:"Transicion JK"
  //: /end
  _GGOR2 #(6) g22 (.I0(w10), .I1(w14), .Z(w7));   //: @(284,232) /sn:0 /w:[ 1 1 0 ]
  //: IN g0 (K) @(37,256) /sn:0 /w:[ 0 ]
  //: comment g12 @(720,56) /sn:0
  //: /line:"Como pone en internet(no funciona)"
  //: /end
  FlipFlopD g18 (.Reloj(Reloj), .D(w7), .W(w12), .nQ(nQ), .Q(Q));   //: @(374, 257) /sz:(129, 78) /sn:0 /p:[ Li0>1 Li1>1 Bi0>1 Ro0<0 Ro1<0 ]
  _GGAND2 #(6) g33 (.I0(!R), .I1(J), .Z(w5));   //: @(106,207) /sn:0 /w:[ 3 0 0 ]
  //: joint g30 (w8) @(645, 239) /w:[ -1 2 12 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin Suma
module Suma(AcarreoE, B, Suma, AcarreoS, A);
//: interface  /sz:(67, 60) /bd:[ Ti0>AcarreoE(33/67) Li0>B(37/60) Li1>A(15/60) Bo0<AcarreoS(33/67) Ro0<Suma(28/60) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(98,198)(220,198){1}
//: {2}(224,198)(254,198){3}
//: {4}(258,198)(374,198){5}
//: {6}(378,198)(408,198){7}
//: {8}(412,198)(438,198){9}
//: {10}(442,198)(475,198)(475,235){11}
//: {12}(440,200)(440,210)(441,210)(441,236){13}
//: {14}(410,200)(410,235){15}
//: {16}(376,200)(376,210)(377,210)(377,235){17}
//: {18}(256,200)(256,210)(254,210)(254,232){19}
//: {20}(222,200)(222,210)(220,210)(220,232){21}
input A;    //: /sn:0 {0}(436,236)(436,136){1}
//: {2}(438,134)(470,134)(470,235){3}
//: {4}(434,134)(406,134){5}
//: {6}(402,134)(370,134){7}
//: {8}(366,134)(282,134){9}
//: {10}(278,134)(215,134){11}
//: {12}(211,134)(103,134){13}
//: {14}(213,136)(213,146)(215,146)(215,232){15}
//: {16}(280,136)(280,146)(284,146)(284,232){17}
//: {18}(368,136)(368,146)(372,146)(372,235){19}
//: {20}(404,136)(404,146)(405,146)(405,235){21}
input AcarreoE;    //: /sn:0 {0}(232,46)(232,110)(246,110){1}
//: {2}(250,110)(288,110){3}
//: {4}(292,110)(378,110){5}
//: {6}(382,110)(414,110){7}
//: {8}(418,110)(444,110){9}
//: {10}(448,110)(480,110)(480,235){11}
//: {12}(446,112)(446,236){13}
//: {14}(416,112)(416,122)(415,122)(415,235){15}
//: {16}(380,112)(380,122)(382,122)(382,235){17}
//: {18}(290,112)(290,122)(289,122)(289,232){19}
//: {20}(248,112)(248,122)(249,122)(249,232){21}
output AcarreoS;    //: /sn:0 {0}(247,433)(247,366)(251,366)(251,351){1}
output Suma;    //: /sn:0 {0}(433,432)(433,359)(428,359)(428,344){1}
wire w14;    //: /sn:0 {0}(425,323)(425,301)(410,301)(410,256){1}
wire w20;    //: /sn:0 {0}(475,256)(475,308)(435,308)(435,323){1}
wire w8;    //: /sn:0 {0}(286,253)(286,320)(256,320)(256,330){1}
wire w17;    //: /sn:0 {0}(430,323)(430,300)(441,300)(441,257){1}
wire w11;    //: /sn:0 {0}(377,256)(377,308)(420,308)(420,323){1}
wire w2;    //: /sn:0 {0}(217,253)(217,321)(246,321)(246,330){1}
wire w5;    //: /sn:0 {0}(251,253)(251,330){1}
//: enddecls

  _GGOR4 #(10) g8 (.I0(w20), .I1(w17), .I2(w14), .I3(w11), .Z(Suma));   //: @(428,334) /sn:0 /R:3 /w:[ 1 0 0 1 1 ]
  _GGAND3 #(8) g4 (.I0(!AcarreoE), .I1(B), .I2(!A), .Z(w14));   //: @(410,246) /sn:0 /R:3 /w:[ 15 15 21 1 ]
  //: IN g13 (AcarreoE) @(232,44) /sn:0 /R:3 /w:[ 0 ]
  _GGAND3 #(8) g3 (.I0(AcarreoE), .I1(!B), .I2(!A), .Z(w11));   //: @(377,246) /sn:0 /R:3 /w:[ 17 17 19 0 ]
  _GGAND2 #(6) g2 (.I0(AcarreoE), .I1(A), .Z(w8));   //: @(286,243) /sn:0 /R:3 /w:[ 19 17 0 ]
  _GGAND2 #(6) g1 (.I0(B), .I1(AcarreoE), .Z(w5));   //: @(251,243) /sn:0 /R:3 /w:[ 19 21 0 ]
  //: joint g16 (AcarreoE) @(248, 110) /w:[ 2 -1 1 20 ]
  //: IN g11 (B) @(96,198) /sn:0 /w:[ 0 ]
  //: joint g28 (AcarreoE) @(446, 110) /w:[ 10 -1 9 12 ]
  //: OUT g10 (Suma) @(433,429) /sn:0 /R:3 /w:[ 0 ]
  //: joint g27 (B) @(440, 198) /w:[ 10 -1 9 12 ]
  //: joint g19 (AcarreoE) @(290, 110) /w:[ 4 -1 3 18 ]
  _GGAND3 #(8) g6 (.I0(AcarreoE), .I1(B), .I2(A), .Z(w20));   //: @(475,246) /sn:0 /R:3 /w:[ 11 11 3 0 ]
  //: OUT g9 (AcarreoS) @(247,430) /sn:0 /R:3 /w:[ 0 ]
  _GGOR3 #(8) g7 (.I0(w8), .I1(w5), .I2(w2), .Z(AcarreoS));   //: @(251,341) /sn:0 /R:3 /w:[ 1 1 1 1 ]
  //: joint g20 (A) @(368, 134) /w:[ 7 -1 8 18 ]
  //: joint g15 (B) @(222, 198) /w:[ 2 -1 1 20 ]
  //: joint g25 (B) @(410, 198) /w:[ 8 -1 7 14 ]
  //: joint g17 (B) @(256, 198) /w:[ 4 -1 3 18 ]
  //: joint g14 (A) @(213, 134) /w:[ 11 -1 12 14 ]
  _GGAND3 #(8) g5 (.I0(!AcarreoE), .I1(!B), .I2(A), .Z(w17));   //: @(441,247) /sn:0 /R:3 /w:[ 13 13 0 1 ]
  //: joint g24 (AcarreoE) @(416, 110) /w:[ 8 -1 7 14 ]
  //: joint g21 (B) @(376, 198) /w:[ 6 -1 5 16 ]
  //: joint g23 (A) @(404, 134) /w:[ 5 -1 6 20 ]
  //: joint g26 (A) @(436, 134) /w:[ 2 -1 4 1 ]
  //: joint g22 (AcarreoE) @(380, 110) /w:[ 6 -1 5 16 ]
  _GGAND2 #(6) g0 (.I0(B), .I1(A), .Z(w2));   //: @(217,243) /sn:0 /R:3 /w:[ 21 15 0 ]
  //: joint g18 (A) @(280, 134) /w:[ 9 -1 10 16 ]
  //: IN g12 (A) @(101,134) /sn:0 /w:[ 13 ]

endmodule
//: /netlistEnd

//: /netlistBegin ALU1bit
module ALU1bit(B, A, C, AcarreoS, AcarreoE, Sa);
//: interface  /sz:(87, 60) /bd:[ Ti0>C[2:0](66/87) Ti1>AcarreoE(31/87) Li0>B(36/60) Li1>A(21/60) Bo0<AcarreoS(32/87) Ro0<Sa(31/60) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(319,334)(276,334)(276,333)(246,333){1}
//: {2}(242,333)(211,333)(211,332)(203,332){3}
//: {4}(201,330)(201,163)(461,163){5}
//: {6}(465,163)(502,163){7}
//: {8}(463,165)(463,182)(503,182){9}
//: {10}(201,334)(201,379)(88,379){11}
//: {12}(244,335)(244,352)(260,352){13}
input A;    //: /sn:0 {0}(420,245)(407,245)(407,160){1}
//: {2}(409,158)(479,158){3}
//: {4}(483,158)(502,158){5}
//: {6}(481,160)(481,177)(503,177){7}
//: {8}(405,158)(186,158)(186,157)(80,157){9}
input AcarreoE;    //: /sn:0 {0}(433,56)(433,214)(454,214)(454,229){1}
output Sa;    //: /sn:0 {0}(716,201)(901,201)(901,199)(916,199){1}
input [2:0] C;    //: /sn:0 {0}(#:694,69)(#:694,35){1}
supply0 w2;    //: /sn:0 {0}(662,207)(593,207){1}
//: {2}(591,205)(591,198)(662,198){3}
//: {4}(589,207)(579,207)(579,217)(662,217){5}
//: {6}(591,209)(591,236){7}
//: {8}(593,238)(662,238){9}
//: {10}(591,240)(591,264){11}
output AcarreoS;    //: /sn:0 {0}(454,291)(454,348)(465,348)(465,363){1}
wire w6;    //: /sn:0 {0}(523,161)(647,161)(647,167)(662,167){1}
wire w7;    //: /sn:0 {0}(524,180)(647,180)(647,179)(662,179){1}
wire w16;    //: /sn:0 {0}(361,341)(406,341)(406,267)(420,267){1}
wire w3;    //: /sn:0 {0}(340,323)(340,120)(682,120){1}
//: {2}(684,118)(684,75){3}
//: {4}(684,122)(684,146)(683,146)(683,159){5}
wire w0;    //: /sn:0 {0}(704,75)(704,144)(705,144)(705,159){1}
wire w1;    //: /sn:0 {0}(694,75)(694,159){1}
wire w8;    //: /sn:0 {0}(662,228)(555,228)(555,230)(545,230){1}
//: {2}(543,228)(543,187)(662,187){3}
//: {4}(543,232)(543,258)(489,258){5}
wire w22;    //: /sn:0 {0}(276,352)(319,352){1}
//: enddecls

  Mux3 g8 (.C2(w3), .C1(w1), .C0(w0), .E7(w2), .E6(w8), .E5(w2), .E4(w2), .E3(w2), .E2(w8), .E1(w7), .E0(w6), .Sal(Sa));   //: @(663, 160) /sz:(52, 85) /sn:0 /p:[ Ti0>5 Ti1>1 Ti2>1 Li0>9 Li1>0 Li2>5 Li3>0 Li4>3 Li5>3 Li6>1 Li7>1 Ro0<0 ]
  //: IN g4 (B) @(86,379) /sn:0 /w:[ 11 ]
  //: joint g13 (w8) @(543, 230) /w:[ 1 2 -1 4 ]
  //: IN g3 (A) @(78,157) /sn:0 /w:[ 9 ]
  //: GROUND g2 (w2) @(591,270) /sn:0 /w:[ 11 ]
  //: IN g1 (C) @(694,33) /sn:0 /R:3 /w:[ 1 ]
  //: joint g16 (A) @(407, 158) /w:[ 2 -1 8 1 ]
  _GGAND2 #(6) g11 (.I0(A), .I1(B), .Z(w6));   //: @(513,161) /sn:0 /w:[ 5 7 0 ]
  Mux1 g10 (.C(w3), .E1(w22), .E0(B), .Sal(w16));   //: @(320, 324) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Li0>1 Li1>0 Ro0<0 ]
  //: joint g19 (B) @(244, 333) /w:[ 1 -1 2 12 ]
  //: OUT g6 (AcarreoS) @(465,360) /sn:0 /R:3 /w:[ 1 ]
  Suma g9 (.AcarreoE(AcarreoE), .A(A), .B(w16), .AcarreoS(AcarreoS), .Suma(w8));   //: @(421, 230) /sz:(67, 60) /sn:0 /p:[ Ti0>1 Li0>0 Li1>1 Bo0<0 Ro0<5 ]
  assign {w3, w1, w0} = C; //: CONCAT g7  @(694,70) /sn:0 /R:1 /w:[ 3 0 0 0 ] /dr:0 /tp:0 /drp:0
  //: joint g20 (w3) @(684, 120) /w:[ -1 2 1 4 ]
  //: joint g15 (B) @(463, 163) /w:[ 6 -1 5 8 ]
  //: joint g17 (B) @(201, 332) /w:[ 3 4 -1 10 ]
  //: joint g14 (A) @(481, 158) /w:[ 4 -1 3 6 ]
  //: IN g5 (AcarreoE) @(433,54) /sn:0 /R:3 /w:[ 0 ]
  //: joint g21 (w2) @(591, 238) /w:[ 8 7 -1 10 ]
  //: joint g22 (w2) @(591, 207) /w:[ 1 2 4 6 ]
  //: OUT g0 (Sa) @(913,199) /sn:0 /w:[ 1 ]
  _GGNBUF #(2) g18 (.I(B), .Z(w22));   //: @(266,352) /sn:0 /w:[ 13 0 ]
  _GGOR2 #(6) g12 (.I0(A), .I1(B), .Z(w7));   //: @(514,180) /sn:0 /w:[ 7 9 0 ]

endmodule
//: /netlistEnd

